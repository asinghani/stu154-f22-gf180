* NGSPICE file created from user_proj.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

.subckt user_proj io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2]
+ io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37]
+ io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0]
+ la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3155_ _0135_ net75 ttA_1.top.data\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout56_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2106_ _0352_ _0354_ _0356_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_3086_ _0066_ net112 ttA_0.data\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1997__C _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _0287_ _0288_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _0893_ _1002_ _1005_ _0924_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3132__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1693__A1 ttA_1.top.backend.rptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3282__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2945__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2531__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1684__A1 ttA_1.top.backend.wptr_gray\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1739__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2936__A1 ttA_0.data\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ _0862_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ _0284_ _0720_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3155__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1606_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2586_ ttA_0.io_out\[6\] _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2164__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout127 net1 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1537_ _1089_ _1090_ _1091_ _1083_ net8 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout105 net107 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3207_ ttA_1.top.backend.wptr_gray1\[3\] _0018_ net29 ttA_1.top.backend.wptr_gray2\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1675__A1 ttA_1.top.frontend.wptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3138_ _0118_ net35 ttA_0.prog\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3069_ _0049_ net69 ttA_1.top.data\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1978__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3019__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2858__I _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3268__294 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2593__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2261__C _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3178__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0585_ _0614_ _0604_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout106_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2768__I _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2371_ _0561_ _0539_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1657__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2909__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2707_ _0517_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2638_ _0402_ _0705_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2569_ _0359_ _0373_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2845__B1 ttA_4.active_duty\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1648__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2346__C _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2588__I _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1887__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1887__B2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1639__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ _1357_ _1460_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2064__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1871_ _1381_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2367__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0585_ _0601_ _0589_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2354_ _1334_ _1396_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2285_ _0496_ _0498_ _0500_ _0495_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2871__I _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _1418_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2781__I _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2972_ _1012_ _1026_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2037__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2714__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_250 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ _1350_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xuser_proj_261 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_272 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_283 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1854_ ttA_4.pwm_signal _1380_ _1381_ ttA_2.io_out\[0\] _1341_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1785_ _1308_ _1314_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ ttA_0.prog\[11\]\[1\] _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2021__I ttA_0.io_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout86_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2956__I _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2337_ _1104_ _1077_ _1370_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2268_ _0485_ _0486_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2276__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2199_ _0438_ _0435_ _0439_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3239__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2503__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2114__S1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1570_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3240_ _0203_ net81 ttA_0.data\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2050__S0 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3171_ _0151_ net105 ttA_0.data\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _0315_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2053_ _0287_ _0305_ _0289_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2258__A1 ttA_0.data\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2955_ _0546_ _0000_ _0945_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1906_ _1340_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2430__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2886_ _0904_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1837_ _1362_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1768_ _1280_ _1299_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ ttA_1.top.backend.wptr_gray2\[2\] _1232_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2619__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3061__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput20 net20 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2032__S0 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2660__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ ttA_0.data\[12\]\[0\] _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2671_ _0816_ _0740_ _0752_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2963__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1622_ _1124_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1553_ net8 _1083_ net5 net4 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3223_ _0186_ net97 ttA_6.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _0134_ net95 ttA_1.top.data\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2105_ _0297_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3085_ _0065_ net107 ttA_0.data\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2036_ _1431_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3084__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2938_ ttA_0.data\[13\]\[1\] _1003_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2954__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2869_ _1088_ _0950_ _0951_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2945__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2259__C _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2723_ _0862_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _0699_ _0721_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1605_ _1081_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2585_ _0374_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1536_ net4 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout117 net125 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout106 net107 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3206_ ttA_1.top.backend.wptr_gray1\[2\] _0017_ net29 ttA_1.top.backend.wptr_gray2\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1675__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3137_ _0117_ net35 ttA_0.prog\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3068_ _0048_ net69 ttA_1.top.data\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2019_ _0263_ _0271_ _1520_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2863__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2615__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3040__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ _1332_ _0376_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2854__B2 ttA_4.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1621__C _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3122__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2909__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2706_ _0328_ _0347_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1593__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2637_ _0733_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3272__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2568_ _0326_ _0473_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _0534_ _0659_ _0661_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2845__B2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2845__A1 ttA_4.active_duty\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1648__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1584__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1722__B _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2109__I _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3145__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1870_ _1342_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1683__I ttA_1.top.frontend.wptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2422_ _0599_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1878__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2353_ _1140_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ ttA_0.data\[8\]\[0\] _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2055__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ ttA_2.io_out\[7\] _1399_ _1472_ _1342_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1566__A1 ttA_2.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2818__A1 ttA_0.data\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3168__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2971_ _1122_ _1014_ _0816_ _1016_ _1025_ _1018_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_251 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_240 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1922_ ttA_6.counter\[1\] _1386_ _1438_ _1351_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_262 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_273 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_284 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_295 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1853_ net11 _1335_ _1336_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1784_ _1272_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _0580_ _0584_ _0587_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout79_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2336_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2267_ _0328_ _0475_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2177__C _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2198_ ttA_1.top.data\[5\]\[1\] _0434_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3271__291 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2368__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__A2 _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2042__I2 ttA_0.prog\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1950__A1 ttA_2.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2050__S1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3170_ _0150_ net103 ttA_0.data\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2121_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2052_ ttA_0.prog\[12\]\[1\] ttA_0.prog\[13\]\[1\] ttA_0.prog\[14\]\[1\] ttA_0.prog\[15\]\[1\]
+ _0298_ _0299_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__2792__I ttA_0.prog\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2954_ _0942_ _0928_ _1013_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1905_ ttA_2.io_out\[3\] _1399_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2885_ _0965_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1836_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1767_ _1294_ _1298_ _1270_ _1272_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__3275__D _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1698_ ttA_1.top.backend.wptr_gray2\[0\] ttA_1.top.backend.rptr_b2g.gray\[0\] _1239_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2319_ ttA_0.data\[6\]\[3\] _0520_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I io_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2032__S1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__A1 ttA_2.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2948__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1956__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2670_ _0741_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1621_ _1144_ _1149_ _1174_ _1126_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ _1100_ _1102_ _1103_ _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3222_ _0185_ _0027_ net44 ttA_1.top.backend.wptr_gray\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3153_ _0133_ net83 ttA_0.prog\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2104_ ttA_0.data\[12\]\[0\] ttA_0.data\[14\]\[0\] ttA_0.data\[13\]\[0\] ttA_0.data\[15\]\[0\]
+ _0330_ _0293_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3084_ _0064_ net111 ttA_0.data\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2035_ ttA_0.prog\[12\]\[0\] ttA_0.prog\[13\]\[0\] ttA_0.prog\[14\]\[0\] ttA_0.prog\[15\]\[0\]
+ _1330_ _1394_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2651__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__I ttA_0.io_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2471__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _0888_ _1002_ _1004_ _0924_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2868_ ttA_0.prog\[2\]\[3\] _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1819_ ttA_6.counter\[7\] _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2799_ _0914_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2167__A1 ttA_0.data\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2646__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2381__B _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1905__A1 ttA_2.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2330__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2633__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2722_ _0848_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2653_ _1500_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2584_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1604_ _1086_ _1156_ _1158_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1535_ net5 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net122 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout107 net110 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3205_ ttA_1.top.backend.wptr_gray1\[1\] _0016_ net28 ttA_1.top.backend.wptr_gray2\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2321__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3136_ _0116_ net35 ttA_0.prog\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3067_ _0047_ net73 ttA_1.top.data\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2018_ ttA_0.prog\[4\]\[2\] ttA_0.prog\[5\]\[2\] ttA_0.prog\[6\]\[2\] ttA_0.prog\[7\]\[2\]
+ _0259_ _1393_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2388__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2615__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3074__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2130__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2303__A1 ttA_0.data\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2705_ _0385_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0755_ _0773_ _0777_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2790__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2567_ _1508_ _1501_ _0391_ _1470_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2040__I _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1896__A3 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2498_ ttA_0.prog\[6\]\[0\] _0660_ _0651_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2975__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3119_ _0099_ net65 ttA_0.prog\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1584__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3193__D ttA_1.top.backend.rptr_b2g.gray\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2885__I _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2772__A1 ttA_0.data\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout111_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2524__A1 ttA_0.prog\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1958__S0 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2352_ _0546_ _0541_ _0547_ _0548_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2795__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ _0497_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1998_ _1248_ _1510_ _1517_ _1340_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2063__I0 ttA_0.data\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2763__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2619_ _0688_ _0704_ _0766_ _0682_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2118__I1 ttA_0.data\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2506__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3112__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1959__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2970_ _1434_ _0641_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xuser_proj_241 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_230 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1921_ _1363_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xuser_proj_252 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_263 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_274 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_285 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_296 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_1852_ _1338_ _1335_ net10 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2993__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1783_ _1309_ _1312_ _1270_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2404_ _0585_ _0586_ _0576_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2335_ _1332_ _1396_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2266_ _0378_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2197_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1869__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2736__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3135__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3285__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2403__I _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2042__I3 ttA_0.prog\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2120_ _0366_ _0368_ _0370_ _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _1417_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2953_ _0593_ _0848_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1904_ _1426_ _1427_ _1367_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2966__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2884_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1835_ _1338_ _1335_ _1336_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__I0 ttA_0.prog\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1766_ _1295_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3158__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2718__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1697_ _1238_ ttA_1.top.backend.rptr_b2g.gray\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout91_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2318_ _0503_ _0519_ _0523_ _0516_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2249_ _0343_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2185__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2024__I3 ttA_0.prog\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput22 net22 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2379__B _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2645__B1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2948__A1 ttA_4.active_duty\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2948__B2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1620__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1620_ _1147_ _1129_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2133__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1551_ net5 _1100_ _1101_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3221_ _0184_ _0026_ net45 ttA_1.top.frontend.wptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_119_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3152_ _0132_ net59 ttA_0.prog\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2103_ _0292_ _0355_ _1432_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3083_ _0063_ net106 ttA_0.data\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2034_ _0263_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2939__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ ttA_0.data\[13\]\[0\] _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2867_ _0955_ _0949_ _0956_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1818_ ttA_6.counter\[11\] _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2798_ _0914_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _1271_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1669__A1 ttA_1.top.frontend.rptr_gray2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2094__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2291__C _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2721_ _0860_ _0852_ _0861_ _0859_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2652_ _0344_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2798__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1603_ ttA_2.io_out\[7\] _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2583_ _0326_ _0473_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1534_ net6 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout119 net122 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3204_ ttA_1.top.backend.wptr_gray1\[0\] _0015_ net31 ttA_1.top.backend.wptr_gray2\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3135_ _0115_ net54 ttA_0.prog\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3066_ _0046_ net74 ttA_1.top.data\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout54_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2017_ _1416_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2482__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2919_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2560__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2379__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2000__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2067__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2704_ _1509_ _0704_ _0828_ _0847_ _0848_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2635_ _0775_ _0757_ _0728_ _1477_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2566_ _0312_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2497_ _0658_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3118_ _0098_ net71 ttA_0.prog\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2991__I _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3049_ _1303_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2533__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2387__B _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2406__I ttA_0.prog\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2221__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2420_ _0581_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout104_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1958__S1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2351_ _0515_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2282_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2288__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1997_ _1250_ _1513_ _1516_ _1231_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2212__A1 ttA_1.top.data\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2063__I1 ttA_0.data\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2763__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _0707_ _0765_ _0704_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2549_ _0280_ _0282_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1890__I ttA_0.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2515__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2118__I2 ttA_0.data\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2279__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3064__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2506__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_242 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_231 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_220 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1920_ _1346_ _1360_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xuser_proj_253 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_264 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_275 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_297 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__2993__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1851_ _1368_ _1371_ _1375_ _1376_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_129_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_286 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ _1292_ _1311_ _1290_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _0583_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2334_ _1140_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2265_ _0349_ _0364_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2196_ _0397_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3087__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2046__I _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2984__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2672__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2035__S0 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2050_ ttA_0.prog\[8\]\[1\] ttA_0.prog\[9\]\[1\] ttA_0.prog\[10\]\[1\] ttA_0.prog\[11\]\[1\]
+ _0298_ _0299_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2952_ _0931_ _0390_ _1009_ _0433_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1903_ _1149_ _1371_ _1409_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _0611_ _0644_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _1357_ _1359_ _1360_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1638__C _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1696_ ttA_1.top.backend.rptr\[1\] ttA_1.top.backend.rptr\[0\] _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2026__S0 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2317_ ttA_0.data\[6\]\[2\] _0520_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2248_ _0448_ _0469_ _0472_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2179_ _1143_ ttA_1.top.frontend.wptr\[0\] _1220_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2957__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3102__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput23 net23 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2893__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2395__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2645__B2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2948__A2 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _1104_ ttA_2.io_out\[0\] _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3220_ _0183_ _0025_ net47 ttA_1.top.frontend.wptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3151_ _0131_ net59 ttA_0.prog\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2102_ ttA_0.data\[8\]\[0\] ttA_0.data\[9\]\[0\] ttA_0.data\[10\]\[0\] ttA_0.data\[11\]\[0\]
+ _0329_ _0330_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3082_ _0062_ net106 ttA_0.data\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2033_ _1417_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3125__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _1001_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2866_ _0592_ _0950_ _0951_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1817_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2797_ _0914_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3275__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1748_ _1270_ _1272_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1679_ ttA_1.top.frontend.wptr\[2\] _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2875__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3052__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1669__A2 ttA_1.top.backend.wptr_gray\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3043__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2720_ ttA_0.data\[14\]\[3\] _0853_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2651_ _0744_ _0760_ _0717_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1983__I _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1602_ _1085_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2582_ _0725_ _0727_ _0729_ _0701_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1533_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3203_ _0175_ net84 ttA_0.data\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3134_ _0114_ net34 ttA_0.prog\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3065_ _0045_ net73 ttA_1.top.data\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2016_ ttA_0.prog\[0\]\[2\] ttA_0.prog\[1\]\[2\] ttA_0.prog\[2\]\[2\] ttA_0.prog\[3\]\[2\]
+ _0266_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout47_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3034__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2918_ _0989_ _0990_ _1401_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1596__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2849_ ttA_4.active_duty\[4\] _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1893__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1977__I3 ttA_1.top.data\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2551__A3 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2067__A2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3016__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ _1377_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2634_ _0701_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2602__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ _0693_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2496_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3117_ _0097_ net92 ttA_0.prog\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3048_ _1062_ _1072_ _1073_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__C _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 net102 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout80 net81 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2422__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1732__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2350_ ttA_0.prog\[15\]\[3\] _0542_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2281_ _0412_ _0476_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2460__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1996_ _1235_ ttA_1.top.data\[2\]\[2\] _1515_ _1233_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2212__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2063__I2 ttA_0.data\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2332__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1971__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0724_ _0730_ _0747_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2548_ _0273_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2479_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2242__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2054__I2 ttA_0.prog\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1962__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_232 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_210 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_221 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_243 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_265 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_254 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_276 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _1377_ _1373_ _1166_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1781_ _1279_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2152__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ _1176_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1705__A1 ttA_1.top.backend.rptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ _0505_ _0527_ _0532_ _0533_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2101__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ _0405_ _0478_ _0483_ _0484_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2195_ _0433_ _0435_ _0436_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2755__C _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1979_ ttA_0.io_out\[6\] _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2062__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1850__B _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2672__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2424__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__S1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2951_ _0932_ _1012_ _1009_ _0549_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1902_ _0003_ _1403_ _1424_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2882_ ttA_0.prog\[1\]\[0\] _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1833_ ttA_6.counter\[11\] _1344_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2179__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1764_ beepboop.inst.counter\[6\] _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1695_ ttA_1.top.backend.wptr_gray2\[1\] ttA_1.top.backend.rptr_b2g.gray\[1\] _1237_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__S1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3054__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout77_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2316_ _0501_ _0519_ _0522_ _0516_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ ttA_1.top.data\[0\]\[2\] _0468_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2103__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2178_ _1197_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput24 net24 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2590__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2520__I _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2581__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2333__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3150_ _0130_ net59 ttA_0.prog\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3081_ _0061_ net46 ttA_1.top.data\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2101_ _0297_ _0353_ _0255_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2032_ ttA_0.prog\[8\]\[0\] ttA_0.prog\[9\]\[0\] ttA_0.prog\[10\]\[0\] ttA_0.prog\[11\]\[0\]
+ _1330_ _1394_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2934_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2865_ ttA_0.prog\[2\]\[2\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1816_ ttA_6.counter\[15\] ttA_6.counter\[14\] ttA_6.counter\[13\] ttA_6.counter\[12\]
+ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_102_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2796_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ _1274_ _1278_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1678_ _1224_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3279_ _0242_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2627__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2315__A1 ttA_0.data\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout127_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2650_ _1477_ _0794_ _0795_ _0770_ _0768_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1601_ _1088_ _1121_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2581_ _0688_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2160__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1532_ _1081_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3202_ _0174_ net82 ttA_0.data\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3133_ _0113_ net36 ttA_0.prog\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3064_ _0044_ net74 ttA_1.top.data\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2015_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3242__CLK net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2917_ _0930_ _0937_ _0934_ _0988_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2793__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2848_ ttA_4.active_duty\[5\] _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2779_ _0582_ _0644_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2784__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2536__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2155__I _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2702_ _0756_ _0836_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2633_ _0391_ _0778_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2564_ _0708_ _0709_ _0710_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2527__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2495_ _0550_ _0657_ _0642_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3116_ _0096_ net71 ttA_0.prog\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3047_ beepboop.inst.counter\[9\] beepboop.inst.counter\[8\] _1070_ _1073_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_110_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3007__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2065__I _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__I0 ttA_0.data\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2766__A1 ttA_0.data\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2518__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3288__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout70 net77 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout92 net94 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout81 net82 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _0385_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2594__B _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1989__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _1478_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2748__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2616_ _0749_ _0755_ _0759_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2547_ _0689_ _0690_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1723__A2 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2920__A1 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2478_ _0641_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2054__I3 ttA_0.prog\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_233 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_200 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_211 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_222 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_244 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_266 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_255 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1650__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_277 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ beepboop.inst.counter\[3\] _1273_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2401_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2332_ _0515_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2263_ _0421_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2194_ ttA_1.top.data\[5\]\[0\] _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1978_ _1248_ _1498_ _1430_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A3 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1880__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2188__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2950_ _0407_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2881_ beepboop.inst.counter\[0\] _0962_ _0963_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1623__A1 ttA_2.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1901_ _1129_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1832_ _1353_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2179__A2 ttA_1.top.frontend.wptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1763_ _1284_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ _1236_ ttA_1.top.backend.rptr_b2g.gray\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ ttA_0.data\[6\]\[1\] _0520_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2246_ _0446_ _0469_ _0471_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2177_ _0405_ _0414_ _0419_ _0422_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__I _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput25 net25 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput14 net14 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2590__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2581__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ _0060_ net67 ttA_1.top.data\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2100_ ttA_0.data\[4\]\[0\] ttA_0.data\[6\]\[0\] ttA_0.data\[5\]\[0\] ttA_0.data\[7\]\[0\]
+ _0330_ _0293_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0273_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2158__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2933_ _0379_ _0850_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2864_ _0953_ _0949_ _0954_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1815_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2795_ _1368_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1746_ beepboop.inst.counter\[1\] beepboop.inst.counter\[0\] _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ ttA_1.top.backend.wptr_gray\[3\] _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3171__CLK net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3278_ _0241_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2229_ _0446_ _0458_ _0460_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2260__A1 ttA_0.data\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2563__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2687__B _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2079__A1 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1610__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2251__A1 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1600_ _1122_ _1139_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _0693_ _0725_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1531_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3291__287 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3201_ _0173_ net83 ttA_0.data\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3132_ _0112_ net33 ttA_0.prog\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3063_ _0043_ net73 ttA_1.top.data\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2014_ ttA_0.io_out\[1\] _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2916_ ttA_4.counter\[5\] ttA_4.counter\[4\] _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2847_ ttA_4.active_duty\[4\] _0929_ ttA_4.active_duty\[3\] _0930_ _0939_ _0940_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2351__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2778_ ttA_0.prog\[3\]\[0\] _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1729_ _1100_ _1079_ _1264_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3067__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2536__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2701_ _0767_ _0841_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2632_ _0696_ _0283_ _0714_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2563_ _1470_ _0359_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2083__S0 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2494_ _1419_ _0256_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3115_ _0095_ net72 ttA_0.prog\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3046_ _1304_ _1070_ _1306_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout52_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2066__I1 ttA_0.data\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2081__I _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2518__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2965__B _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2206__A1 ttA_1.top.data\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout71 net76 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout60 net62 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout82 net85 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2693__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1938__C _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1994_ ttA_1.top.data\[3\]\[2\] _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2115__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2615_ _0762_ _0711_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2056__S0 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _0689_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2920__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3165__RN _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2684__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3029_ _1276_ _1059_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2436__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2076__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2804__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3105__CLK net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__S0 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2675__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2427__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_201 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_212 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_223 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_245 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_234 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_267 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_256 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1650__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_278 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2400_ _0581_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout102_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ ttA_0.data\[4\]\[3\] _0528_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2262_ ttA_0.data\[9\]\[3\] _0479_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2193_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2666__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3128__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1977_ ttA_1.top.data\[4\]\[1\] ttA_1.top.data\[5\]\[1\] ttA_1.top.data\[6\]\[1\]
+ ttA_1.top.data\[7\]\[1\] _1481_ _1479_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__3278__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ _0420_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2657__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1699__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2896__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2880_ net13 _1281_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1900_ _1406_ _1407_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1623__A2 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2820__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _1351_ _1348_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2179__A3 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ _1291_ _1293_ _1276_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_129_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1693_ ttA_1.top.backend.rptr\[2\] ttA_1.top.backend.rptr\[1\] _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2314_ _0496_ _0519_ _0521_ _0516_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ ttA_1.top.data\[0\]\[1\] _0468_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2176_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2811__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2575__B1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput15 net15 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2878__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2529__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2102__I0 ttA_0.data\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2030__A2 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2869__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2030_ _1433_ _0276_ _0278_ _0280_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2932_ _0992_ _1000_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2863_ _0632_ _0950_ _0951_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1814_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2794_ _0911_ _0902_ _0912_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2902__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _1275_ beepboop.inst.counter\[4\] _1276_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__B _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1676_ _1208_ _1209_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout82_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3277_ _0240_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2228_ ttA_1.top.data\[2\]\[1\] _0457_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2088__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2159_ _0381_ _0405_ _0406_ _0408_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3037__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2812__I _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2012__A2 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2079__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2722__I _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _1080_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3200_ _0172_ net81 ttA_0.data\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3131_ _0111_ net64 ttA_0.prog\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3062_ _0042_ net68 ttA_1.top.data\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2013_ ttA_0.io_out\[0\] _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2915_ _0988_ _0928_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2846_ _0931_ ttA_4.counter\[3\] _0932_ ttA_4.counter\[2\] _0936_ _0938_ _0939_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2777_ _0898_ _0890_ _0899_ _0897_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1728_ _1079_ _1260_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1659_ ttA_1.top.frontend.wptr\[1\] _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2807__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1992__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2472__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3161__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0842_ _0843_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2631_ _0733_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2562_ _1500_ _0343_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2083__S1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ _0655_ _0646_ _0656_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3114_ _0094_ net92 ttA_0.prog\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3045_ _1067_ _1071_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout45_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1974__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2829_ _0915_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net79 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout72 net76 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1965__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout94 net96 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1717__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2142__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2447__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2445__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _1252_ ttA_1.top.data\[0\]\[2\] _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0689_ _0719_ _0692_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2056__S1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1526__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2381__A1 ttA_0.prog\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0690_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3057__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2476_ _1434_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2684__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3028_ _1301_ _1057_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2436__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2092__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2047__S1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2124__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2675__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_202 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_213 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_224 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_246 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_235 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_257 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_268 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_279 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A1 ttA_6.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2330_ _0503_ _0527_ _0531_ _0525_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2261_ _0400_ _0478_ _0482_ _0422_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2192_ _1208_ _1228_ _1222_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2666__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3213__D net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1976_ _1250_ _1493_ _1496_ ttA_1.top.backend.rptr\[2\] _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1944__A4 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2528_ ttA_0.prog\[4\]\[3\] _0676_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _0585_ _0629_ _0617_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3222__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2648__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ ttA_6.counter\[3\] _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1761_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1692_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3208__D ttA_1.top.backend.wptr_gray\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2313_ ttA_0.data\[6\]\[0\] _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1804__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2244_ _0442_ _0469_ _0470_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2175_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3245__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2811__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1959_ _1234_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2575__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput27 net27 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput16 net16 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2878__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1714__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1550__A2 ttA_2.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2102__I1 ttA_0.data\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2280__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2318__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3118__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3268__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2931_ ttA_4.counter\[5\] _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2862_ ttA_0.prog\[2\]\[1\] _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1813_ _1337_ _1339_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2190__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2404__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2793_ _0623_ _0903_ _0905_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1744_ beepboop.inst.counter\[7\] beepboop.inst.counter\[6\] _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1675_ ttA_1.top.frontend.wptr\[0\] _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2309__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1534__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3276_ _0239_ _0032_ net65 ttA_2.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _0442_ _0458_ _0459_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2158_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2089_ _0289_ _0332_ _0337_ _0339_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2720__A1 ttA_0.data\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2087__I0 ttA_0.data\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2787__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1762__A2 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__I0 ttA_0.prog\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3090__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ _0110_ net41 ttA_0.prog\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2711__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3061_ _0041_ net68 ttA_1.top.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2012_ _0263_ _0264_ _1431_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__I0 ttA_0.data\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2914_ ttA_4.counter\[0\] _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2845_ ttA_4.active_duty\[2\] _0937_ ttA_4.active_duty\[1\] _0934_ _0938_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2776_ ttA_0.data\[10\]\[3\] _0891_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1727_ _1190_ _1261_ _1262_ _1084_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1658_ ttA_1.top.frontend.wptr\[2\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2702__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1589_ ttA_2.io_out\[5\] _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3259_ _0222_ net119 ttA_6.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2823__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2769__A1 ttA_0.data\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout125_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _0756_ _0774_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2561_ ttA_0.io_out\[7\] _0326_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2492_ _0623_ _0648_ _0651_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3113_ _0093_ net92 ttA_0.prog\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3044_ _1304_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ _0926_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ _0857_ _0880_ _0884_ _0886_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1726__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2151__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2981__C _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__A1 ttA_1.top.frontend.wptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout40 net49 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout73 net75 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout62 net63 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout51 net52 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1653__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2463__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ _1481_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1807__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2613_ _0745_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2544_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2381__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2475_ _0537_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3027_ _0962_ _1058_ _1059_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3151__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2548__I _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1883__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_203 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_214 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2283__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_247 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_236 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_225 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_269 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_258 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1938__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2060__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ ttA_0.data\[9\]\[2\] _0479_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2191_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2666__A3 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2193__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1975_ _1252_ _1494_ _1495_ _1479_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2354__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0437_ _0675_ _0679_ _0548_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2458_ _0627_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2389_ _0554_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1617__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2290__A1 ttA_0.data\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2831__I _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1640__I1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2345__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1553__B1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2278__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2281__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ beepboop.inst.counter\[4\] _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3197__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1691_ ttA_1.top.backend.rptr\[0\] _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2312_ _0518_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ ttA_1.top.data\[0\]\[0\] _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2174_ _1372_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1820__I ttA_6.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2272__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1958_ ttA_1.top.data\[4\]\[0\] ttA_1.top.data\[5\]\[0\] ttA_1.top.data\[6\]\[0\]
+ ttA_1.top.data\[7\]\[0\] _1478_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1889_ _1376_ _1375_ _1405_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput17 net17 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1838__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1730__I ttA_2.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2102__I2 ttA_0.data\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2510__B _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2930_ ttA_4.counter\[4\] _0996_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2861_ _0947_ _0949_ _0952_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1812_ _1338_ net9 _1336_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2792_ ttA_0.prog\[3\]\[3\] _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1743_ beepboop.inst.counter\[3\] _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1674_ _1142_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3275_ _0238_ _0031_ net64 ttA_2.io_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_100_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ ttA_1.top.data\[2\]\[0\] _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout68_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2157_ _1377_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2088_ _0333_ _0340_ _0289_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2556__I _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2236__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2087__I1 ttA_0.data\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__B _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3235__CLK net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ _0040_ net108 ttA_0.data\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2011_ ttA_0.prog\[12\]\[2\] ttA_0.prog\[13\]\[2\] ttA_0.prog\[14\]\[2\] ttA_0.prog\[15\]\[2\]
+ _0259_ _1393_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2227__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0986_ _0978_ _0987_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2844_ ttA_4.counter\[2\] _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2775_ _0404_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1726_ _1133_ _1130_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1657_ _1098_ _1086_ _1204_ _1207_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ _0221_ net121 ttA_6.counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2376__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ ttA_1.top.data\[4\]\[1\] _0443_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3189_ ttA_1.top.frontend.rptr_gray1\[1\] _0004_ net38 ttA_1.top.frontend.rptr_gray2\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__A1 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3258__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2286__I _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__S0 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout118_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2560_ _1476_ _0374_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2491_ ttA_0.prog\[7\]\[3\] _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2696__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3112_ _0092_ net71 ttA_0.prog\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2196__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3043_ _1062_ _1069_ _1070_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2448__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _0926_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2758_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1709_ _1248_ _1245_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2923__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2689_ _0831_ _0832_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2687__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__A2 ttA_1.top.frontend.wptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout30 net31 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout41 net44 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2611__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout63 net78 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout52 net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout96 net101 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout85 net91 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__B2 ttA_4.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ ttA_1.top.data\[1\]\[2\] _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2612_ _0311_ _0691_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _1433_ _0296_ _0301_ _0286_ _0290_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ _0318_ _0535_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1823__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2669__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout50_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3026_ beepboop.inst.counter\[2\] _1057_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2829__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_204 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_215 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_248 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_237 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_226 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_259 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2513__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2899__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2190_ _1197_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1974_ _1235_ ttA_1.top.data\[0\]\[1\] _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1818__I ttA_6.counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2051__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ ttA_0.prog\[4\]\[2\] _0676_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2457_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2388_ _0549_ _0572_ _0574_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2114__I0 ttA_0.data\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _0960_ _1050_ _1051_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1617__A2 ttA_2.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2814__A1 ttA_0.data\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1553__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1553__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2294__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2281__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2033__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ ttA_1.top.backend.rptr\[1\] _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1792__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1544__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2311_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3291_ net287 clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2173_ ttA_0.data\[0\]\[3\] _0415_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1976__C ttA_1.top.backend.rptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1957_ ttA_1.top.backend.rptr\[1\] _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1888_ _1362_ _1392_ _1414_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3291__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2509_ _0666_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2971__B1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2289__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3164__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2860_ _0647_ _0950_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1811_ _1338_ net10 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2791_ _0909_ _0902_ _0910_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ beepboop.inst.counter\[5\] _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3274_ _0237_ _0030_ net43 ttA_2.io_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_113_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2225_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2156_ ttA_0.data\[1\]\[3\] _0387_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2087_ ttA_0.data\[12\]\[2\] ttA_0.data\[14\]\[2\] ttA_0.data\[13\]\[2\] ttA_0.data\[15\]\[2\]
+ _0334_ _0335_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__2245__A2 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2989_ _1385_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_135_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__B _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3187__CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1995__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__I2 ttA_0.prog\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2172__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2010_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2078__I2 ttA_0.data\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2912_ _1088_ _0979_ _0980_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1986__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1986__B2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2843_ ttA_4.active_duty\[1\] _0934_ ttA_4.active_duty\[0\] _0935_ _0936_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2774_ _0895_ _0890_ _0896_ _0897_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ _1131_ _1106_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1656_ _1138_ _1206_ _1157_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1587_ _1104_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2163__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout80_I net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3257_ _0220_ net99 ttA_6.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _0397_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3188_ ttA_1.top.frontend.rptr_gray1\[0\] _0003_ net45 ttA_1.top.frontend.rptr_gray2\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2466__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2139_ _1476_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__I2 ttA_0.data\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1729__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2154__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2209__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1968__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3202__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__S1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__A1 ttA_0.prog\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ _0653_ _0646_ _0654_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2696__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3111_ _0091_ net72 ttA_0.prog\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3042_ _1284_ beepboop.inst.counter\[6\] _1065_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2145__C _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2826_ _0926_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2384__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _0420_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1708_ _1231_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2688_ _1500_ _0374_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1639_ _1122_ _1187_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1990__S0 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__3225__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout64 net70 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout42 net44 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout53 net56 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net99 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2611__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout86 net89 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2375__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2127__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2678__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2297__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2850__A2 ttA_4.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ ttA_1.top.data\[4\]\[2\] ttA_1.top.data\[5\]\[2\] ttA_1.top.data\[6\]\[2\]
+ ttA_1.top.data\[7\]\[2\] _1478_ _1479_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_127_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2611_ _0756_ _0757_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2366__A1 ttA_0.prog\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2542_ _0311_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2473_ ttA_0.prog\[7\]\[0\] _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2669__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3025_ _1273_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2935__I _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout43_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2670__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ _0917_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1580__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_205 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_238 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_216 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_227 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_249 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2596__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2060__A3 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2348__A1 _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1924__I ttA_6.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ ttA_1.top.data\[1\]\[1\] _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2339__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2525_ _0432_ _0675_ _0678_ _0548_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_115_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2456_ _0581_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3070__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ ttA_0.prog\[12\]\[0\] _0573_ _0566_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2511__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3008_ ttA_6.counter\[8\] _1049_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2114__I1 ttA_0.data\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2578__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2333__C _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2502__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2569__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3093__CLK net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3290_ net288 clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1544__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2310_ _0487_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2741__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2241_ _0424_ _0462_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0400_ _0414_ _0418_ _0408_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2434__B _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1956_ _1234_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2104__S0 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1887_ _1396_ _1397_ _1399_ _1130_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput19 net19 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2508_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2439_ _0612_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2971__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1810_ net11 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2790_ _0620_ _0903_ _0905_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1672_ _1214_ _1216_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2962__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2714__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3273_ _0236_ _0029_ net64 ttA_2.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2224_ _0456_ _0424_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2155_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2086_ _0292_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2988_ _1034_ _1035_ _1037_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_107_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1939_ _1347_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2953__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1995__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1747__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2944__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3131__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3281__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ ttA_0.prog\[0\]\[3\] _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2842_ ttA_4.counter\[0\] _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2773_ _0885_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1724_ _1164_ _1198_ _1132_ _1256_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1655_ _1180_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2003__I _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1586_ ttA_2.io_out\[4\] _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout73_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3256_ _0219_ net90 ttA_0.data\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2207_ _0442_ _0444_ _0445_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3187_ _0167_ net37 ttA_0.prog\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1998__B _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _0381_ _0386_ _0388_ _0390_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2069_ ttA_0.data\[0\]\[3\] ttA_0.data\[1\]\[3\] ttA_0.data\[2\]\[3\] ttA_0.data\[3\]\[3\]
+ _1330_ _1394_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2069__I3 ttA_0.data\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1729__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3154__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2145__A2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3110_ _0090_ net92 ttA_0.prog\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3041_ _1297_ _1065_ _1295_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1656__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2825_ _0926_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3177__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2756_ ttA_0.data\[15\]\[2\] _0881_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1707_ _1247_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2687_ _0687_ _0751_ _0343_ _1476_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1638_ _1164_ _1188_ _1189_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1572__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1569_ _1090_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1895__B2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1895__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__S1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3239_ _0202_ net82 ttA_0.data\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout32 net2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout65 net70 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout54 net56 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout76 net77 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout87 net89 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__C _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2375__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2127__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2610_ _0687_ _0361_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2366__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ _0273_ _0283_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2472_ _0638_ _0628_ _0639_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1877__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3024_ _1279_ _0962_ _1057_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1629__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout36_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2808_ _0917_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0871_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__I _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3022__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2293__A1 ttA_0.data\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_206 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_239 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_217 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_228 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2284__A1 ttA_0.data\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2771__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1972_ ttA_1.top.data\[2\]\[1\] ttA_1.top.data\[3\]\[1\] _1481_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2704__C _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2339__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2524_ ttA_0.prog\[4\]\[1\] _0676_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2455_ _1419_ _0570_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2386_ _0571_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2511__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3007_ _1436_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2114__I2 ttA_0.data\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2578__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3017__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2502__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2569__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2240_ _0448_ _0464_ _0467_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2171_ ttA_0.data\[0\]\[2\] _0415_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1955_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__3249__D _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2104__S1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2006__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1886_ _1400_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2507_ _0561_ _0657_ _0642_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2438_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2369_ _0440_ _0552_ _0560_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2248__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__C _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2098__S0 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3060__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1740_ beepboop.inst.counter\[2\] _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1671_ _1212_ ttA_1.top.backend.wptr_gray\[1\] _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3272_ _0235_ _0028_ net66 ttA_2.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ _1208_ _1228_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2478__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__S0 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2154_ _0402_ _0382_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ ttA_0.data\[8\]\[2\] ttA_0.data\[9\]\[2\] ttA_0.data\[10\]\[2\] ttA_0.data\[11\]\[2\]
+ _0329_ _0294_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2650__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2987_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1938_ ttA_6.counter\[4\] _1438_ _1349_ _1350_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2953__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1869_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2641__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1747__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2910_ _0984_ _0978_ _0985_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2841_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2772_ ttA_0.data\[10\]\[2\] _0891_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1723_ _1167_ _1080_ _1259_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1654_ _1163_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1585_ _1133_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2699__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3255_ _0218_ net87 ttA_0.data\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2206_ ttA_1.top.data\[4\]\[0\] _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout66_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3186_ _0166_ net53 ttA_0.prog\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1674__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2068_ ttA_0.data\[4\]\[3\] ttA_0.data\[6\]\[3\] ttA_0.data\[5\]\[3\] ttA_0.data\[7\]\[3\]
+ _1395_ _1331_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2623__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2903__B _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3040_ _1067_ _1068_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2853__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2605__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2824_ _0915_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__I ttA_0.io_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2755_ _0855_ _0880_ _0883_ _0877_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ _1232_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2686_ _0804_ _0806_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1637_ _1081_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1568_ _1089_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3238_ _0201_ net119 ttA_4.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3169_ _0149_ net89 ttA_0.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout44 net48 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2633__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout33 net34 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout66 net68 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2352__C _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1958__I0 ttA_1.top.data\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1583__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2859__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3271__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2527__C _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3012__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2540_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2471_ _0623_ _0629_ _0634_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3023_ beepboop.inst.counter\[1\] beepboop.inst.counter\[0\] _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2009__I ttA_0.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout29_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2807_ _0915_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2738_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2669_ _0809_ _0706_ _0738_ _0810_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2817__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_229 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_207 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_218 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2596__A3 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__C _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3167__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1971_ _1477_ _1343_ _1489_ _1492_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2523_ _0534_ _0675_ _0677_ _0548_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2454_ ttA_0.prog\[8\]\[0\] _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2385_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3006_ _0960_ _1048_ _1049_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1578__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2027__A2 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _0395_ _0414_ _0417_ _0408_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2782__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ ttA_0.io_out\[5\] _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1885_ _1401_ _1402_ _1405_ _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout96_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _0430_ _0659_ _0665_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1940__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2437_ _0581_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2368_ ttA_0.prog\[14\]\[3\] _0553_ _0557_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2299_ ttA_0.data\[5\]\[0\] _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2248__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2906__B _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1972__S _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__B2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2088__B _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1998__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2107__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2098__S1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ ttA_1.top.backend.wptr_gray\[3\] ttA_1.top.frontend.rptr_gray2\[3\] _1217_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3271_ net291 net124 ttA_6.counter\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _1514_ _0451_ _0455_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2022__S1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2153_ _1159_ _0383_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _0333_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2986_ ttA_6.counter\[1\] ttA_6.counter\[0\] _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1937_ _1351_ _1348_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1868_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1799_ beepboop.inst.counter\[11\] _1270_ _1282_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_131_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1913__A1 ttA_6.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2469__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3228__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2641__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2880__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2840_ ttA_4.counter\[1\] _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2632__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2396__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2771_ _0399_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1722_ _1255_ _1258_ _1080_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _1160_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2148__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__B _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1584_ _1123_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3254_ _0217_ net87 ttA_0.data\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3185_ _0165_ net53 ttA_0.prog\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2136_ _1372_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2067_ _0318_ _0319_ _1434_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1586__I ttA_2.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2969_ _1022_ _1024_ _1012_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__A1 ttA_0.prog\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2366__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2917__A3 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2550__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2302__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2853__A2 ttA_4.pwm_signal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2823_ _0917_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2369__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2754_ ttA_0.data\[15\]\[1\] _0881_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1705_ ttA_1.top.backend.rptr\[2\] _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ _1471_ _0741_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1636_ _1165_ _1132_ _1163_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3273__D _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ _1087_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2541__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3237_ _0200_ net119 ttA_4.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3168_ _0148_ net88 ttA_0.data\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2119_ _0333_ _0371_ _0255_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3099_ _0079_ net114 ttA_0.data\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout45 net47 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout34 net36 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout56 net63 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout78 net79 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2205__I _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1583__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2096__B _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2599__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2470_ ttA_0.prog\[8\]\[3\] _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2523__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3022_ _1056_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2806_ _0916_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1864__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2737_ _0412_ _0850_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2668_ _0811_ _0812_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1619_ _1165_ _1170_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2599_ _1509_ _0732_ _0743_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2514__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2909__B _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_208 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_219 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2753__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1970_ _1397_ _1454_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2116__S0 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2992__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ ttA_0.prog\[4\]\[0\] _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2744__A1 ttA_0.data\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0622_ _0613_ _0624_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2384_ _0570_ _0539_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3005_ ttA_6.counter\[7\] _1046_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout41_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2983__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2035__I0 ttA_0.prog\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2735__A1 ttA_0.data\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__I3 ttA_0.prog\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2374__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3270__292 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_139_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1701__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3284__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1679__I ttA_1.top.frontend.wptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _1469_ _1475_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1884_ _1403_ _1406_ _1407_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1628__B _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ ttA_0.prog\[6\]\[3\] _0660_ _0662_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2436_ _1420_ _0561_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ _0438_ _0552_ _0559_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2298_ _0508_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3157__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1998__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2947__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2123__I _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ net292 net123 ttA_6.counter\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1922__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _1196_ _0450_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1686__A1 ttA_1.top.frontend.wptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _1508_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2083_ ttA_0.data\[4\]\[2\] ttA_0.data\[6\]\[2\] ttA_0.data\[5\]\[2\] ttA_0.data\[7\]\[2\]
+ _0334_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2635__B1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2985_ _0959_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2938__A1 ttA_0.data\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1936_ _1387_ _1456_ _1457_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_135_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1867_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1798_ _1293_ _1318_ _1277_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _1420_ _0550_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1677__A1 ttA_1.top.backend.wptr_gray\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2208__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1601__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2093__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2632__A3 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2770_ _0893_ _0890_ _0894_ _0886_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1721_ _1164_ _1173_ _1256_ _1257_ _1122_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _1099_ _1112_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ _1126_ _1132_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3253_ _0216_ net86 ttA_0.data\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _1225_ _1228_ _0424_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3184_ _0164_ net53 ttA_0.prog\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2135_ ttA_0.data\[1\]\[0\] _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2066_ ttA_0.data\[12\]\[3\] ttA_0.data\[14\]\[3\] ttA_0.data\[13\]\[3\] ttA_0.data\[15\]\[3\]
+ _1395_ _1331_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2623__A3 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1867__I _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2968_ _0809_ _1016_ _1023_ _1018_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1919_ _1435_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2899_ _0626_ _0643_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2075__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2917__A4 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2401__I _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__A1 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2550__A2 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2822_ _0898_ _0919_ _0925_ _0924_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2369__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2753_ _0849_ _0880_ _0882_ _0877_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1704_ _1233_ _1235_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1636__B _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2684_ _0775_ _0758_ _0807_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1635_ _1136_ _1146_ _1133_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ ttA_2.io_out\[7\] _1094_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2311__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2541__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout71_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3236_ _0199_ net121 ttA_4.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3167_ _0147_ _0002_ net73 ttA_2.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3098_ _0078_ net114 ttA_0.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2118_ ttA_0.data\[4\]\[1\] ttA_0.data\[6\]\[1\] ttA_0.data\[5\]\[1\] ttA_0.data\[7\]\[1\]
+ _0274_ _0335_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ _1433_ _0296_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2057__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout46 net47 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout35 net36 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout68 net70 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout79 net127 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout57 net62 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_136_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1958__I2 ttA_1.top.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1546__B net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2377__B _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2296__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2220__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3021_ _1056_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2287__A1 ttA_0.data\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2306__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2805_ _0916_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2736_ _0860_ _0864_ _0870_ _0869_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2667_ _1501_ _0809_ _0779_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1618_ _1124_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2041__I _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2598_ _0745_ _0720_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2514__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1549_ _1091_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3219_ _0182_ _0024_ net41 ttA_1.top.frontend.wptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_209 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2216__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2202__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2886__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2554__C _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2116__S1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3063__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2992__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2521_ _0674_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2452_ _0623_ _0614_ _0617_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2052__S0 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2383_ _1334_ _0376_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3004_ _1387_ _1046_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout34_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ _0404_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2499__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2671__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3086__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1952_ _1243_ _1430_ _1397_ _1471_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1883_ _1168_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2504_ _0428_ _0659_ _0664_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2435_ ttA_0.prog\[9\]\[0\] _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2366_ ttA_0.prog\[14\]\[2\] _0553_ _0557_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2297_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2016__S0 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__A2 ttA_1.top.backend.rptr_b2g.gray\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2947__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3101__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2007__S0 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _0438_ _0451_ _0454_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2279__C _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1686__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2883__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2151_ _0381_ _0400_ _0401_ _0390_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2082_ _0258_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2635__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2635__B2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2984_ ttA_6.counter\[1\] _1386_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1935_ _1456_ _1447_ _1387_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1866_ ttA_0.io_out\[1\] _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1797_ _1308_ _1322_ _1323_ _1325_ _1314_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2418_ ttA_0.prog\[10\]\[0\] _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1677__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _1180_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2626__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3124__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2843__B ttA_4.active_duty\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _1167_ _1109_ _1107_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1141_ _1086_ _1195_ _1202_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1582_ _1133_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ _0215_ net93 ttA_0.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1922__B _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ _1197_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2856__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3183_ _0163_ net80 ttA_0.data\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _0380_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2065_ _0287_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2084__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3033__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2967_ _0318_ _0536_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1918_ _1436_ _1440_ _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1595__A1 ttA_2.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2898_ ttA_0.prog\[0\]\[0\] _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ _1372_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2075__A2 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3024__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__I _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2821_ ttA_0.data\[2\]\[3\] _0920_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2752_ ttA_0.data\[15\]\[0\] _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1703_ _1125_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2799__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2683_ _0801_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1634_ _1185_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1565_ _1095_ _1096_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_141_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3235_ _0198_ net122 ttA_4.counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3166_ _0146_ _0001_ net74 ttA_2.io_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout64_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3097_ _0077_ net113 ttA_0.data\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2039__I ttA_0.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2117_ _0257_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2057__A2 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ _0297_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout36 net37 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3006__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net62 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2296__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2393__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2048__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2412__I _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1731__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3020_ _1056_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1798__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2804_ _0916_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2735_ ttA_0.data\[3\]\[3\] _0865_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2666_ _1502_ _0809_ _0757_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ _1143_ ttA_2.io_out\[0\] _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2597_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1548_ _1090_ _1101_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3218_ _0181_ net51 ttA_0.prog\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3149_ _0129_ net60 ttA_0.prog\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1961__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2441__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout114_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1952__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1952__B2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2451_ _1087_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1981__I _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ _0440_ _0563_ _0569_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2052__S1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ _1039_ _1046_ _1047_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2718_ _0857_ _0852_ _0858_ _0859_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2987__I _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2649_ _0751_ _0769_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2671__B _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2026__I2 ttA_0.prog\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2137__I _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _1425_ _1400_ _1408_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1882_ _1373_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2503_ ttA_0.prog\[6\]\[2\] _0660_ _0662_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2600__I _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2434_ _0608_ _0600_ _0609_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _0433_ _0552_ _0558_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2296_ _0379_ _0487_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2653__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__A1 ttA_0.data\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1916__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2016__S1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3053__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2007__S1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2150_ ttA_0.data\[1\]\[2\] _0387_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ _0267_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2635__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _0898_ _1028_ _1033_ _0823_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1934_ _1456_ _1448_ _1358_ ttA_6.counter\[2\] _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2399__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1865_ _1364_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1796_ _1316_ _1324_ _1315_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3076__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout94_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2417_ _0595_ _0584_ _0596_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2348_ _0437_ _0541_ _0545_ _0533_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2486__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2279_ _0405_ _0489_ _0494_ _0495_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2626__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2314__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2415__I ttA_0.prog\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3099__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1650_ _1196_ _1201_ _1157_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1581_ _1098_ _1128_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3251_ _0214_ net93 ttA_0.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2305__A1 ttA_0.data\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _0440_ _0435_ _0441_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3182_ _0162_ net80 ttA_0.data\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2133_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2064_ _1418_ _0316_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2753__C _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2966_ _0593_ _1014_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_190 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1917_ ttA_6.counter\[9\] _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2897_ _0974_ _0966_ _0975_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1848_ _1142_ _1076_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1595__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1779_ beepboop.inst.counter\[10\] beepboop.inst.counter\[9\] _1277_ _1309_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_137_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3241__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__A1 ttA_1.top.data\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0895_ _0919_ _0923_ _0924_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2751_ _0879_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1702_ _1237_ _1239_ _1240_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1577__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2682_ _0709_ _0825_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2774__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1633_ _1115_ _1096_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2526__A1 ttA_0.prog\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1564_ ttA_2.io_out\[6\] _1094_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3234_ _0197_ net118 ttA_4.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2748__C _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3165_ _0145_ _0000_ net94 ttA_2.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3096_ _0076_ net113 ttA_0.data\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2116_ ttA_0.data\[0\]\[1\] ttA_0.data\[1\]\[1\] ttA_0.data\[2\]\[1\] ttA_0.data\[3\]\[1\]
+ _1329_ _0334_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_fanout57_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3264__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2047_ ttA_0.prog\[4\]\[0\] ttA_0.prog\[5\]\[0\] ttA_0.prog\[6\]\[0\] ttA_0.prog\[7\]\[0\]
+ _0298_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout37 net50 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout59 net61 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2949_ _1011_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1894__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2056__I0 ttA_0.prog\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1559__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3287__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2995__A1 ttA_6.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2803_ _0916_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2747__A1 ttA_0.data\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _0857_ _0864_ _0868_ _0869_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2665_ _0735_ _0728_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1616_ _1166_ _1167_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2596_ _0273_ _0697_ _0698_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_141_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1547_ _1090_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3217_ _0180_ net51 ttA_0.prog\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3148_ _0128_ net55 ttA_0.prog\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3079_ _0059_ net46 ttA_1.top.data\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2977__A1 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2729__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1952__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2450_ ttA_0.prog\[9\]\[3\] _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1704__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ ttA_0.prog\[13\]\[3\] _0564_ _0566_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[14] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3002_ _1456_ _1044_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2968__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2761__C _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ _0681_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1943__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ _0751_ _0769_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2489__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2579_ _0720_ _0715_ _0726_ _0714_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2959__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__I3 ttA_0.prog\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ ttA_2.io_out\[4\] _1398_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1881_ _1406_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2502_ _0423_ _0659_ _0663_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2433_ _1196_ _0601_ _0604_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1689__A1 ttA_1.top.backend.rptr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2364_ ttA_0.prog\[14\]\[1\] _0553_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2350__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2295_ _0505_ _0498_ _0506_ _0507_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2080_ _0262_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2096__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2982_ ttA_0.data\[11\]\[3\] _1029_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1933_ ttA_6.counter\[6\] _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2399__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1864_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1795_ _1292_ _1301_ _1296_ _1291_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2416_ _1196_ _0586_ _0589_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout87_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2347_ ttA_0.prog\[15\]\[2\] _0542_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2278_ _0421_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1834__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__I _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2562__A2 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3170__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2250__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1580_ _1128_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2553__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3250_ _0213_ net93 ttA_0.io_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ ttA_1.top.data\[5\]\[2\] _0434_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3181_ _0161_ net80 ttA_0.data\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2132_ _1471_ _0382_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ ttA_0.data\[8\]\[3\] ttA_0.data\[9\]\[3\] ttA_0.data\[10\]\[3\] ttA_0.data\[11\]\[3\]
+ _1331_ _1395_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_180 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2965_ _1020_ _1021_ _0928_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xuser_proj_191 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1916_ _1357_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2896_ _1088_ _0967_ _0968_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1847_ _1374_ _1371_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1778_ _1302_ _1305_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__I1 ttA_0.data\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2535__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3066__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2471__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2750_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ ttA_1.top.backend.wptr_gray2\[2\] _1232_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2681_ _0344_ _0717_ _0800_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1632_ _1117_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1563_ _1097_ _1114_ _1115_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_126_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3233_ _0196_ net118 ttA_4.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3164_ _0144_ net88 ttA_0.data\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2115_ _0333_ _0367_ _1432_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3095_ _0075_ net113 ttA_0.data\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2046_ _0274_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout38 net40 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3006__A3 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2948_ ttA_4.active_duty\[1\] _0823_ _1009_ _1425_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2879_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2517__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3089__CLK net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A3 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2692__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2802_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2733_ _0681_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2664_ _0778_ _0746_ _0732_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1615_ _1168_ _1130_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2595_ _0733_ _0738_ _0742_ _0731_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1546_ net8 _1082_ net4 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2759__C _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3231__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3216_ _0179_ net51 ttA_0.prog\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2683__A1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ _0127_ net55 ttA_0.prog\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3078_ _0058_ net66 ttA_1.top.data\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2029_ _0263_ _0281_ _1431_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3104__CLK net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2729__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0438_ _0563_ _0568_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3001_ ttA_6.counter\[6\] _1044_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput6 io_in[15] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2665__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1712__I0 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2716_ ttA_0.data\[14\]\[2\] _0853_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2647_ _0767_ _0792_ _0793_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2028__S0 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2578_ _0687_ _0362_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1529_ _1081_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2656__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2408__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3127__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3277__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1880_ net3 _1369_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ ttA_0.prog\[6\]\[1\] _0660_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2432_ ttA_0.prog\[10\]\[3\] _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1689__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2363_ _0555_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ _0421_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2638__A1 _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2877__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2629__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2096__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1843__A2 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3045__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2981_ _0895_ _1028_ _1032_ _0823_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1932_ _1429_ _1455_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1863_ _1385_ ttA_6.counter\[1\] _1386_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1794_ _1291_ _1293_ _1295_ _1297_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2415_ ttA_0.prog\[11\]\[3\] _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__C _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2346_ _0432_ _0541_ _0544_ _0533_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2277_ ttA_0.data\[7\]\[3\] _0490_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2802__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2693__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2712__I _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2200_ _1160_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3180_ _0160_ net80 ttA_0.data\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2131_ _1126_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2062_ _0313_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2964_ _1205_ _1014_ _0784_ _1016_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_181 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_170 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1915_ _1348_ _1438_ _1350_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xuser_proj_192 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2895_ ttA_0.prog\[1\]\[3\] _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _1372_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1777_ _1303_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3290__288 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2329_ ttA_0.data\[4\]\[2\] _0528_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input12_I io_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__A1 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__I _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2083__I2 ttA_0.data\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2223__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1700_ ttA_1.top.backend.rptr\[3\] ttA_1.top.backend.wptr_gray2\[3\] _1241_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2680_ _0796_ _0799_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1982__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1631_ _1097_ _1114_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1562_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3232_ _0195_ net58 ttA_0.prog\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _0143_ net104 ttA_0.data\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ ttA_0.data\[12\]\[1\] ttA_0.data\[14\]\[1\] ttA_0.data\[13\]\[1\] ttA_0.data\[15\]\[1\]
+ _0268_ _0335_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3094_ _0074_ net113 ttA_0.data\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1521__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2045_ _1329_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout28 net30 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout39 net40 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3160__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2947_ _0003_ _1009_ _1010_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2878_ net12 _1288_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_136_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1829_ ttA_6.counter\[7\] _1349_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2453__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1964__A1 _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1606__I _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2141__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2692__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2995__A3 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _1368_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2732_ ttA_0.data\[3\]\[2\] _0865_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2663_ _0473_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2900__I _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1614_ _1127_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2594_ _0739_ _0740_ _0741_ _0733_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1545_ ttA_2.io_out\[1\] _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2380__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3215_ _0178_ net51 ttA_0.prog\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2132__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout62_I net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ _0126_ net60 ttA_0.prog\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3077_ _0057_ net67 ttA_1.top.data\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2028_ ttA_0.prog\[12\]\[3\] ttA_0.prog\[13\]\[3\] ttA_0.prog\[14\]\[3\] ttA_0.prog\[15\]\[3\]
+ _0266_ _0268_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2199__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2810__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3056__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2371__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2362__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput7 io_in[16] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3000_ _1039_ _1044_ _1045_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2665__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2715_ _0399_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ _0392_ _0767_ _0670_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2028__S1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2577_ _0696_ _0283_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1528_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2105__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__I _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3129_ _0109_ net33 ttA_0.prog\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2805__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2540__I _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2344__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2715__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2583__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout112_I net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ _0633_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2431_ _0606_ _0600_ _0607_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2335__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2362_ _0549_ _0552_ _0556_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2293_ ttA_0.data\[8\]\[3\] _0499_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2360__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2574__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2629_ _0775_ _0758_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2326__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2629__A2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3244__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2270__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2317__A1 ttA_0.data\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1614__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2980_ ttA_0.data\[11\]\[2\] _1029_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1931_ _1220_ _1430_ _1343_ _1434_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_128_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1862_ _1359_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 io_in[19] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1793_ _1306_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__S0 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2308__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2414_ _0591_ _0584_ _0594_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2345_ ttA_0.prog\[15\]\[1\] _0542_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2276_ _0400_ _0489_ _0493_ _0484_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3267__CLK net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2090__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2538__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2130_ _0350_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2061_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2175__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3211__D ttA_1.top.backend.wptr_gray\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_160 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2963_ _0570_ _0536_ _1018_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_182 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_171 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1914_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2777__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_proj_193 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2894_ _0972_ _0966_ _0973_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1845_ net95 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ beepboop.inst.counter\[9\] _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout92_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2701__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2328_ _0501_ _0527_ _0530_ _0525_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2259_ _0395_ _0478_ _0481_ _0422_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2813__I _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2969__B _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2723__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2759__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _1086_ _1182_ _1183_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2931__A1 ttA_4.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1734__A2 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1561_ ttA_2.io_out\[4\] _1093_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3231_ _0194_ net57 ttA_0.prog\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3162_ _0142_ net104 ttA_0.data\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ _0257_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1802__I _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3093_ _0073_ net116 ttA_0.data\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2119__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2044_ _0262_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout29 net30 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1670__A1 ttA_1.top.backend.wptr_gray\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2946_ ttA_4.active_duty\[0\] _0000_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2877_ _0003_ _1422_ _0960_ _1386_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1828_ _1345_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1759_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2808__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2150__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2989__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__A3 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2800_ _0914_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2047__I3 ttA_0.prog\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0855_ _0864_ _0867_ _0859_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2662_ _0776_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1613_ _1134_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2593_ _0325_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1544_ _1098_ _1092_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2380__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3214_ _0177_ net97 ttA_4.pwm_signal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3145_ _0125_ net60 ttA_0.prog\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3076_ _0056_ net66 ttA_1.top.data\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2027_ _1416_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2363__I _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2929_ _0992_ _0998_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2362__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3150__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[17] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1625__A1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0855_ _0852_ _0856_ _0682_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1527__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2645_ _0772_ _0783_ _0791_ _0701_ _0784_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2576_ _0697_ _0698_ _0713_ _0723_ _0696_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1527_ net7 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2105__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3128_ _0108_ net33 ttA_0.prog\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3059_ _0039_ net103 ttA_0.data\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1616__A1 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2592__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1552__B1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1855__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2583__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0593_ _0601_ _0604_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout105_I net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__B _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2335__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ ttA_0.prog\[14\]\[0\] _0553_ _0000_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2292_ _0404_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2178__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2099__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3196__CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2628_ ttA_0.io_out\[5\] _0373_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2559_ _0705_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__B _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2262__A1 ttA_0.data\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2565__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _1443_ _1445_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2253__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1861_ _1387_ _1349_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput11 io_in[20] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1792_ _1278_ _1315_ _1320_ _1304_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_128_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2100__S1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3462_ net27 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2413_ _0593_ _0586_ _0589_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1805__I _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2344_ _0534_ _0541_ _0543_ _0533_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2275_ ttA_0.data\[7\]\[2\] _0490_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2492__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2244__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2538__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2060_ _1091_ _1504_ _0284_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2474__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_150 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2962_ _1012_ _1019_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_161 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_183 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_172 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1913_ ttA_6.counter\[3\] ttA_6.counter\[2\] _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2191__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2893_ _0592_ _0967_ _0968_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xuser_proj_194 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1844_ net32 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1775_ _1303_ _1304_ _1295_ _1296_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2085__S0 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1535__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3234__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout85_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ ttA_0.data\[4\]\[1\] _0528_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2258_ ttA_0.data\[9\]\[1\] _0479_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2189_ _0430_ _0426_ _0431_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2465__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2068__I1 ttA_0.data\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3107__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3257__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1560_ ttA_2.io_out\[5\] _1093_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__I0 ttA_1.top.data\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3230_ _0193_ net58 ttA_0.prog\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3161_ _0141_ net88 ttA_0.data\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ ttA_0.data\[8\]\[1\] ttA_0.data\[9\]\[1\] ttA_0.data\[10\]\[1\] ttA_0.data\[11\]\[1\]
+ _1329_ _0334_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3092_ _0072_ net111 ttA_0.data\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2043_ _0292_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2945_ _1266_ _1256_ _0389_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_128_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2876_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1827_ _1346_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1758_ _1275_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1689_ ttA_1.top.backend.rptr\[3\] _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2989__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2824__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2610__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A2 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2601__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ ttA_0.data\[3\]\[1\] _0865_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2661_ _0804_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1612_ _1128_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2592_ _0391_ _0409_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ ttA_2.io_out\[3\] _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2904__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3213_ net3 _0023_ net74 ttA_2.state vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3144_ _0124_ net55 ttA_0.prog\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3075_ _0055_ net45 ttA_1.top.data\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2026_ ttA_0.prog\[8\]\[3\] ttA_0.prog\[9\]\[3\] ttA_0.prog\[10\]\[3\] ttA_0.prog\[11\]\[3\]
+ _0266_ _0268_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0929_ _0996_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2859_ _0904_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2503__B _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[18] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1625__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2822__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1928__A3 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2713_ ttA_0.data\[14\]\[1\] _0853_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2644_ _0746_ _0732_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2575_ _0714_ _0718_ _0712_ _0720_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ net8 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1561__A1 ttA_2.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1543__I ttA_2.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ _0107_ net64 ttA_0.prog\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3058_ _0038_ net108 ttA_0.data\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2009_ ttA_0.io_out\[2\] _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2104__I0 ttA_0.data\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2360_ _0555_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2291_ _0503_ _0498_ _0504_ _0495_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3048__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__C _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1538__I _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A2 _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2627_ _0688_ _0752_ _0740_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2558_ _0695_ _0700_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2489_ _0620_ _0648_ _0651_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2832__I _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2053__B _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3140__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3290__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2253__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1860_ ttA_6.counter\[7\] _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput12 io_in[30] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1791_ _1316_ _1319_ _1277_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2961__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2961__C2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2412_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2343_ ttA_0.prog\[15\]\[0\] _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2274_ _0395_ _0489_ _0492_ _0484_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout30_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2244__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2952__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__A1 ttA_0.data\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1641__I _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3186__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_151 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_140 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2961_ _1198_ _1014_ _0736_ _1016_ _1018_ _1334_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_184 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_173 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_162 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1912_ ttA_6.counter\[8\] _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2892_ ttA_0.prog\[1\]\[2\] _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xuser_proj_195 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1843_ _1370_ net95 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1774_ beepboop.inst.counter\[8\] _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__S1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2162__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout78_I net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2326_ _0496_ _0527_ _0529_ _0525_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2257_ _0386_ _0478_ _0480_ _0422_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2188_ ttA_1.top.data\[6\]\[2\] _0425_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2465__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2068__I2 ttA_0.data\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3059__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2153__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2557__I _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2456__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2292__I _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1967__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2392__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2144__A1 ttA_0.data\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3160_ _0140_ net118 ttA_0.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ _0350_ _0362_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3091_ _0071_ net111 ttA_0.data\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ ttA_0.prog\[0\]\[0\] ttA_0.prog\[1\]\[0\] ttA_0.prog\[2\]\[0\] ttA_0.prog\[3\]\[0\]
+ _0293_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2944_ _0898_ _1002_ _1008_ _1007_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2875_ _1401_ _1345_ _1355_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1826_ _1347_ _1352_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3201__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1757_ _1281_ _1289_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2383__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1688_ ttA_1.top.backend.rptr\[2\] _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _0349_ _0411_ _0375_ _0377_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3289_ net289 clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input10_I io_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2610__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1972__I1 ttA_1.top.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2126__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3224__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0775_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2750__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ _1124_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2591_ _1471_ _0362_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2365__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1542_ ttA_2.io_out\[4\] _1092_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3212_ _0176_ net93 ttA_0.lastdata3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2117__A1 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2197__I _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _0123_ net54 ttA_0.prog\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3074_ _0054_ net66 ttA_1.top.data\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2025_ _0262_ _0277_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _0991_ _0996_ _0997_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2858_ _0948_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1809_ _1335_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2789_ ttA_0.prog\[3\]\[2\] _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2659__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2835__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3247__CLK net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__I _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _0394_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2643_ _0784_ _0786_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2338__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2574_ _0716_ _0717_ _0721_ _0715_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1525_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3126_ _0106_ net33 ttA_0.prog\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout60_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3057_ _0037_ net103 ttA_0.data\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2008_ _0257_ _0260_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2568__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__I _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__S0 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1644__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__A1 ttA_0.data\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ ttA_0.data\[8\]\[2\] _0499_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2475__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2559__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2424__B _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2626_ _0392_ _0705_ _0758_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2557_ _0362_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3092__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2731__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2488_ ttA_0.prog\[7\]\[2\] _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3109_ _0089_ net84 ttA_0.prog\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2098__I0 ttA_0.data\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2970__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput13 io_in[31] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1790_ _1290_ beepboop.inst.counter\[4\] _1318_ _1296_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2961__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout110_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ net7 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2342_ _0540_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2713__A1 ttA_0.data\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2273_ ttA_0.data\[7\]\[1\] _0490_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2138__C _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1549__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1988_ ttA_0.io_out\[7\] _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2952__B2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2609_ _0721_ _0725_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2704__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_141 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_130 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_2960_ _1425_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xuser_proj_152 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_174 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_163 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1911_ ttA_6.counter\[10\] _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2891_ _0970_ _0966_ _0971_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_185 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1842_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_196 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1773_ beepboop.inst.counter\[10\] _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2702__B _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2162__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2325_ ttA_0.data\[4\]\[0\] _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3130__CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2256_ ttA_0.data\[9\]\[0\] _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2187_ _1180_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2663__I _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3280__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1900__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2916__A1 ttA_4.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1719__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3153__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2144__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2110_ _1332_ _0345_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3090_ _0070_ net111 ttA_0.data\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2041_ _0267_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2943_ ttA_0.data\[13\]\[3\] _1003_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2874_ _0913_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1825_ ttA_6.counter\[10\] ttA_6.counter\[9\] ttA_6.counter\[8\] _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1756_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2151__C _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ _1230_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout90_I net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2135__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2308_ _0505_ _0509_ _0514_ _0516_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3288_ net290 clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2239_ ttA_1.top.data\[1\]\[2\] _0463_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1949__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2071__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2374__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3176__CLK net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1885__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2517__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1610_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2590_ _0735_ _0736_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2365__A2 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1541_ ttA_2.io_out\[5\] _1093_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3211_ ttA_1.top.backend.wptr_gray\[3\] _0022_ net28 ttA_1.top.backend.wptr_gray1\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3142_ _0122_ net60 ttA_0.prog\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3073_ _0053_ net45 ttA_1.top.data\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1628__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ ttA_0.prog\[4\]\[3\] ttA_0.prog\[5\]\[3\] ttA_0.prog\[6\]\[3\] ttA_0.prog\[7\]\[3\]
+ _0266_ _0274_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3199__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2926_ ttA_4.counter\[3\] _0994_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2053__A1 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2857_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1808_ net10 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2788_ _0907_ _0902_ _0908_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1739_ beepboop.inst.counter\[11\] _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2347__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2298__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0849_ _0852_ _0854_ _0682_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2642_ _0787_ _0788_ _0748_ _0778_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2573_ _0690_ _0692_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2338__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _1078_ ttA_2.state _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2001__I ttA_0.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3125_ _0105_ net42 ttA_0.prog\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2510__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3056_ _0036_ net108 ttA_0.data\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout53_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2007_ ttA_0.prog\[8\]\[2\] ttA_0.prog\[9\]\[2\] ttA_0.prog\[10\]\[2\] ttA_0.prog\[11\]\[2\]
+ _0259_ _1393_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2274__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2577__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2909_ _0592_ _0979_ _0980_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2067__B _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2104__I2 ttA_0.data\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2265__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2568__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__S1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2256__A1 ttA_0.data\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__A1 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__I ttA_0.prog\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2559__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2625_ _0768_ _0770_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2556_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2487_ _0650_ _0646_ _0652_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3108_ _0088_ net61 ttA_0.prog\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3039_ _1297_ _1065_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2970__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2238__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2410_ ttA_0.prog\[11\]\[2\] _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout103_I net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2341_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2272_ _0386_ _0489_ _0491_ _0484_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2229__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1987_ _1497_ _1499_ _1507_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2952__A2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2608_ _0694_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2704__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2539_ ttA_0.io_out\[4\] _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2468__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2640__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3020__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3188__RN _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_142 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_131 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_153 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_175 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_164 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1910_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2890_ _1205_ _0967_ _0968_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_186 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1841_ net32 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_197 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1772_ _1292_ _1301_ _1290_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2698__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2324_ _0526_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2255_ _0477_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2186_ _0428_ _0426_ _0429_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2916__A2 ttA_4.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0259_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2764__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__A2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2942_ _0895_ _1002_ _1006_ _1007_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0913_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ _1348_ ttA_6.counter\[3\] _1349_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1755_ _1282_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2907__A2 _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2004__I ttA_0.io_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1591__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ ttA_1.top.frontend.wptr\[0\] _1221_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout83_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3287_ _0250_ clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2307_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2238_ _0446_ _0464_ _0466_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2843__A1 ttA_4.active_duty\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ ttA_0.data\[0\]\[1\] _0415_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1885__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2834__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1540_ ttA_2.io_out\[6\] _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3270__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3210_ ttA_1.top.backend.wptr_gray\[2\] _0021_ net28 ttA_1.top.backend.wptr_gray1\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3141_ _0121_ net35 ttA_0.prog\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ _0052_ net43 ttA_1.top.data\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2023_ _1416_ _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2925_ ttA_4.counter\[3\] _0994_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2053__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2856_ _0598_ _0644_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ net9 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2787_ _0632_ _0903_ _0905_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ beepboop.inst.counter\[15\] beepboop.inst.counter\[14\] beepboop.inst.counter\[13\]
+ beepboop.inst.counter\[12\] _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_102_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ ttA_1.top.frontend.rptr_gray2\[0\] ttA_1.top.backend.wptr_gray\[0\] _1216_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1573__I _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2618__B _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2116__I0 ttA_0.data\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2816__A1 ttA_0.data\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3143__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1658__I ttA_1.top.frontend.wptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2710_ ttA_0.data\[14\]\[0\] _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ _1502_ _0736_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1546__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2572_ _0719_ _0692_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1523_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3124_ _0104_ net41 ttA_0.prog\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3055_ _0035_ net103 ttA_0.data\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3166__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _0258_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout46_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2908_ ttA_0.prog\[0\]\[2\] _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2839_ ttA_4.active_duty\[2\] _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1537__B2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2862__I ttA_0.prog\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2017__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1700__A1 ttA_1.top.backend.rptr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2964__B1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2624_ _0768_ _0770_ _0762_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _1402_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2486_ _0632_ _0648_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3107_ _0087_ net59 ttA_0.prog\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2247__A2 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3038_ _0961_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2098__I2 ttA_0.data\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2183__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3018__I _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2022__I2 ttA_0.prog\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1930__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2857__I _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1997__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2525__C _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ _0536_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1921__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ ttA_0.data\[7\]\[0\] _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3204__CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1986_ _1502_ _1342_ _1398_ _1147_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2607_ _0752_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2538_ _0546_ _0683_ _0686_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2677__I _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2469_ _0636_ _0628_ _0637_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3269__293 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2468__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2626__B _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2640__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2361__B _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1903__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2459__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_132 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_154 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_143 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_165 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_176 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1840_ _1076_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xuser_proj_187 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_198 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _1276_ _1273_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2395__A1 ttA_0.prog\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2147__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2698__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2323_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2254_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2185_ ttA_1.top.data\[6\]\[1\] _0425_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2622__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _1367_ _1411_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1576__I _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2310__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2613__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2301__A1 ttA_0.data\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2852__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2941_ _0885_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2780__I _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2872_ _0913_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1823_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ beepboop.inst.counter\[11\] _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _1228_ _1221_ _1229_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1591__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout76_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3286_ _0249_ clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2306_ _0420_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ ttA_1.top.data\[1\]\[1\] _0463_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2843__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2168_ _0386_ _0414_ _0416_ _0408_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2099_ _0292_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2531__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2834__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2598__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2770__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3140_ _0120_ net54 ttA_0.prog\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2775__I _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3071_ _0051_ net42 ttA_1.top.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ ttA_0.prog\[0\]\[3\] ttA_0.prog\[1\]\[3\] ttA_0.prog\[2\]\[3\] ttA_0.prog\[3\]\[3\]
+ _0258_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2589__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2924_ _0992_ _0994_ _0995_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2855_ ttA_0.prog\[2\]\[0\] _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1806_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2015__I _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2786_ ttA_0.prog\[3\]\[1\] _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1737_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2761__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1668_ _1215_ ttA_1.top.backend.wptr_gray\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1599_ _1140_ _1146_ _1151_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ net293 net123 ttA_6.counter\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2116__I1 ttA_0.data\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2052__I0 ttA_0.prog\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2504__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1794__A2 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout126_I net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0392_ _0705_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2571_ _0690_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1522_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2743__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3123_ _0103_ net42 ttA_0.prog\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3054_ _0034_ net108 ttA_0.data\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2005_ ttA_0.io_out\[0\] _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2907_ _0982_ _0978_ _0983_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2838_ ttA_4.active_duty\[3\] _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2769_ ttA_0.data\[10\]\[1\] _0891_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2734__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2348__C _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2364__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2725__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2964__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2623_ _1477_ _0750_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2554_ _0291_ _0302_ _0694_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2716__A1 ttA_0.data\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2192__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2485_ _0633_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3133__CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3106_ _0086_ net83 ttA_0.prog\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3283__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3037_ _1062_ _1065_ _1066_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2098__I3 ttA_0.data\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2955__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2912__B _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2707__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2022__I3 ttA_0.prog\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2946__A1 ttA_4.active_duty\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3156__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2270_ _0488_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2783__I _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1985_ _1409_ _1505_ _1400_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2937__A1 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2606_ _0753_ _0731_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2537_ ttA_1.top.data\[7\]\[2\] _1223_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2468_ _0620_ _0629_ _0634_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2399_ _1420_ _0536_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2642__B _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1600__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3179__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2156__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2868__I ttA_0.prog\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1667__A1 ttA_1.top.frontend.wptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_133 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_155 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_144 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_166 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_177 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_188 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_199 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ _1300_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2778__I ttA_0.prog\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2322_ _0412_ _0487_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2253_ _0379_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2184_ _0397_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ _1144_ _1398_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1899_ _1078_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2138__A2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2846__B1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1649__A1 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2310__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2377__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ ttA_0.data\[13\]\[2\] _1003_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2871_ _0927_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ ttA_6.counter\[5\] _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2368__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1753_ _1269_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ ttA_1.top.backend.wptr_gray\[0\] _1221_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3285_ _0248_ clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2305_ ttA_0.data\[5\]\[3\] _0510_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2236_ _0442_ _0464_ _0465_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2167_ ttA_0.data\[0\]\[0\] _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2098_ ttA_0.data\[0\]\[0\] ttA_0.data\[1\]\[0\] ttA_0.data\[2\]\[0\] ttA_0.data\[3\]\[0\]
+ _0329_ _0294_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2211__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2295__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2121__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3070_ _0050_ net42 ttA_1.top.data\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ ttA_0.io_out\[1\] _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2589__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2923_ ttA_4.counter\[1\] _0988_ ttA_4.counter\[2\] _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2854_ _0940_ _0944_ _0945_ ttA_4.counter\[5\] _0946_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1805_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2785_ _0900_ _0902_ _0906_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2210__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1736_ beepboop.inst.counter\[10\] beepboop.inst.counter\[9\] beepboop.inst.counter\[8\]
+ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1667_ ttA_1.top.frontend.wptr\[1\] ttA_1.top.frontend.wptr\[0\] _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1598_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2513__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3268_ net294 net123 ttA_6.counter\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3199_ _0171_ _0014_ net31 ttA_1.top.backend.rptr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2219_ ttA_1.top.data\[3\]\[1\] _0450_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2116__I2 ttA_0.data\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2876__I _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2504__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ _0715_ _0716_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1521_ net3 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2786__I ttA_0.prog\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3122_ _0102_ net41 ttA_0.prog\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3053_ _0033_ net90 ttA_0.data\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2259__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2004_ ttA_0.io_out\[2\] _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3062__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _1205_ _0979_ _0980_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2837_ ttA_4.counter\[3\] _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2768_ _0394_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1537__A3 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1719_ _1087_ net7 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2699_ _0688_ _0732_ _0753_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2734__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2042__S0 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2489__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3085__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2413__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2622_ _0745_ _0760_ _0360_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2553_ _0695_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2484_ ttA_0.prog\[7\]\[1\] _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__S0 _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3105_ _0085_ net110 ttA_0.data\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3036_ _1291_ _1063_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2465__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2955__A2 _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2643__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2946__A2 _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1685__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _1403_ _1503_ _1404_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2605_ _0714_ _0745_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3100__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2536_ _0437_ _0683_ _0685_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2467_ ttA_0.prog\[8\]\[2\] _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2398_ _0538_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2974__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _1056_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2642__C _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3050__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2884__I _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A2 ttA_1.top.frontend.wptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_156 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_134 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_145 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_167 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_178 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_189 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3123__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3273__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout101_I net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _0505_ _0519_ _0524_ _0525_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _0328_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2183_ _0423_ _0426_ _0427_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _1248_ _1480_ _1488_ _1430_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1898_ _1367_ _1415_ _1421_ _1423_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ _0570_ _0657_ _0642_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2918__B _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1649__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3146__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2074__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1732__B _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1812__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2870_ _0957_ _0949_ _0958_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1821_ ttA_6.counter\[6\] _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3014__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ beepboop.inst.counter\[6\] _1275_ _1283_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ ttA_1.top.frontend.wptr\[1\] _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__I ttA_0.prog\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1879__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3284_ _0247_ clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2304_ _0503_ _0509_ _0513_ _0507_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ ttA_1.top.data\[1\]\[0\] _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2166_ _0413_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3169__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2097_ _0315_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1868__I _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2999_ _1447_ _1042_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1558__A1 ttA_2.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2402__I _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _0261_ _0265_ _0270_ _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1688__I ttA_1.top.backend.rptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2922_ _0937_ _0933_ _0935_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2853_ _0407_ ttA_4.pwm_signal _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1804_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2784_ _0647_ _0903_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1735_ _1232_ ttA_1.top.backend.rptr_b2g.gray\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2312__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1666_ ttA_1.top.frontend.rptr_gray2\[2\] ttA_1.top.backend.wptr_gray\[2\] _1213_
+ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1597_ _1089_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2468__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout81_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1721__B2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3267_ _0230_ net96 ttA_6.counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3198_ _0170_ _0013_ net30 ttA_1.top.backend.rptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2218_ _1485_ _0451_ _0453_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2116__I3 ttA_0.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2149_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2201__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1703__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3121_ _0101_ net71 ttA_0.prog\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3052_ _1067_ _1075_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2003_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2307__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2431__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2905_ ttA_0.prog\[0\]\[1\] _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2836_ ttA_4.counter\[4\] _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2195__A1 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2767_ _0888_ _0890_ _0892_ _0886_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1718_ _1084_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2698_ _0752_ _0716_ _0785_ _0788_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1649_ _1197_ _1198_ _1171_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2498__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__S1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2973__A3 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2186__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3195__D ttA_1.top.backend.rptr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2110__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2621_ _1470_ _0361_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2177__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2552_ _0693_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1915__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2797__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0640_ _0646_ _0649_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2024__S1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3104_ _0084_ net115 ttA_0.data\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3035_ beepboop.inst.counter\[5\] _1063_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2101__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout44_I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1876__I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2168__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _0885_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2340__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2656__B _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2391__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2285__C _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1983_ _1407_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2604_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2535_ ttA_1.top.data\[7\]\[1\] _1223_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2570__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2320__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2466_ _0631_ _0628_ _0635_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2397_ ttA_0.prog\[11\]\[0\] _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2322__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3018_ _0848_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1600__A3 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2313__A1 ttA_0.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_157 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_146 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_135 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_179 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_168 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2140__I _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ _0515_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2251_ _0314_ _0473_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2304__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2182_ ttA_1.top.data\[6\]\[0\] _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ _1250_ _1484_ _1487_ _1231_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1897_ _1356_ _1422_ _1364_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3098__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1977__S0 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0430_ _0667_ _0673_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2985__I _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2449_ _0619_ _0613_ _0621_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1649__A3 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2534__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1820_ ttA_6.counter\[4\] _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3240__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1751_ beepboop.inst.counter\[7\] _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1682_ _1227_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2525__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2303_ ttA_0.data\[5\]\[2\] _0510_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3283_ _0246_ clknet_1_1__leaf_wb_clk_i beepboop.inst.counter\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2096_ _1127_ _1407_ _0314_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__I _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ ttA_6.counter\[5\] _1042_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1949_ _1078_ _1401_ _1373_ _1400_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2516__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3263__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1558__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2755__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2118__S0 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ _0992_ _0993_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2852_ ttA_4.active_duty\[5\] _0555_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1803_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2783_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1734_ _1265_ _1080_ _1268_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2746__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1665_ ttA_1.top.frontend.rptr_gray2\[2\] ttA_1.top.backend.wptr_gray\[2\] ttA_1.top.backend.wptr_gray\[1\]
+ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1596_ _1126_ _1148_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ _0229_ net98 ttA_6.counter\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout74_I net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _0452_ _0451_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3197_ _0169_ _0012_ net31 ttA_1.top.backend.rptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__3286__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2148_ _1502_ _0382_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2079_ _0257_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2737__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2268__A3 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__I0 ttA_0.prog\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2728__A1 ttA_0.data\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3159__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1703__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _0100_ net65 ttA_0.prog\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2288__C _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3051_ _1303_ _1073_ beepboop.inst.counter\[11\] _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2002_ _1520_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2967__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2904_ _0976_ _0978_ _0981_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _0862_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1648__B _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2766_ ttA_0.data\[10\]\[0\] _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1717_ _1153_ _1134_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2697_ _0784_ _0716_ _0773_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1942__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1648_ _1176_ _1178_ _1153_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1579_ ttA_2.io_out\[2\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3249_ _0212_ net83 ttA_0.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2958__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1621__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ _0703_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2143__I _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2016__I3 ttA_0.prog\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2551_ _0696_ _0697_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2482_ _0647_ _0648_ _0634_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3103_ _0083_ net112 ttA_0.data\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3034_ _1062_ _1063_ _1064_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2746__C _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2101__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout37_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2818_ ttA_0.data\[2\]\[2\] _0920_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2749_ _0485_ _0486_ _0850_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1915__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1851__B2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1851__A1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__A1 ttA_2.io_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2159__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1982_ _1149_ _1377_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2534_ _0432_ _0683_ _0684_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2570__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2465_ _0632_ _0629_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2396_ _0430_ _0572_ _0579_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2322__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3017_ _0862_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2086__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1833__A1 ttA_6.counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2492__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2561__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2667__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_147 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_136 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_169 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_158 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2250_ _0318_ _0345_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1965_ _1235_ ttA_1.top.data\[2\]\[0\] _1486_ _1233_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2240__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1896_ _1360_ _1361_ _1390_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_134_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__S1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2517_ ttA_0.prog\[5\]\[3\] _0668_ _0670_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2448_ _0620_ _0614_ _0617_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2379_ ttA_0.prog\[13\]\[2\] _0564_ _0566_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2231__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3192__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2534__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1750_ beepboop.inst.counter\[4\] beepboop.inst.counter\[3\] _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2222__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _1225_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2302_ _0501_ _0509_ _0512_ _0507_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3282_ _0245_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2233_ _1222_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2164_ _0348_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2095_ _0328_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3065__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2213__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2997_ _1039_ _1042_ _1043_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1948_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ _1077_ net32 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2061__I _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2516__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2945__B _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2452__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__S0 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3289__289 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3088__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2574__C _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2118__S1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2920_ _0934_ _0988_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2851_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1802_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2782_ _0554_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ _1266_ _1256_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1664_ ttA_1.top.frontend.rptr_gray2\[1\] _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1595_ ttA_2.io_out\[7\] _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2054__S0 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3265_ _0228_ net98 ttA_6.counter\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1721__A3 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _1123_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3196_ _0168_ _0011_ net30 ttA_1.top.backend.rptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2147_ _0397_ _0383_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2078_ ttA_0.data\[0\]\[2\] ttA_0.data\[1\]\[2\] ttA_0.data\[2\]\[2\] ttA_0.data\[3\]\[2\]
+ _0329_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2737__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2673__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1779__A3 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__I1 ttA_0.prog\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3050_ _1067_ _1074_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2001_ ttA_0.io_out\[3\] _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2664__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2416__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2967__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _1198_ _0979_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2834_ _0440_ _0928_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3103__CLK net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2765_ _0889_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1716_ _1253_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2696_ _0816_ _0706_ _0786_ _0810_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1647_ _1140_ _1170_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3253__CLK net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ _1125_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3248_ _0211_ net97 ttA_4.active_duty\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2655__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3179_ _0159_ net86 ttA_0.data\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__S0 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2646__A1 _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3126__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1621__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout117_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2550_ _1432_ _0276_ _0278_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0645_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3102_ _0082_ net112 ttA_0.data\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3033_ _1293_ _1060_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2817_ _0893_ _0919_ _0922_ _0897_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2748_ _0860_ _0872_ _0878_ _0877_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2679_ _1501_ _0798_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_120_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3149__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__A1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2582__C _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1981_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ _0373_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2533_ ttA_1.top.data\[7\]\[0\] _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2103__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2464_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2395_ ttA_0.prog\[12\]\[3\] _0573_ _0576_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1530__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3016_ _1035_ _1055_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1833__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout120 net121 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_134_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1824__A2 ttA_6.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_148 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_137 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_proj_159 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ _1225_ _1209_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2149__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1964_ _1478_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1895_ _1420_ _1397_ _1399_ _1134_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout97_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _0428_ _0667_ _0672_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2447_ net7 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2378_ _0433_ _0563_ _0567_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2432__I ttA_0.prog\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1680_ _1209_ _1222_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1733__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2301_ ttA_0.data\[5\]\[1\] _0510_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3281_ _0244_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ _1208_ _1209_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2163_ _0349_ _0411_ _0378_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2094_ _0314_ _0344_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2996_ _1448_ _1040_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2770__C _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1947_ ttA_0.io_out\[4\] _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1878_ _1403_ _1376_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2498__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1715__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2063__S1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2850_ _0941_ ttA_4.counter\[5\] _0942_ ttA_4.counter\[4\] _0389_ _0943_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1801_ ttA_0.io_out\[0\] _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2781_ _0901_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1732_ _1079_ _1131_ _1171_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1663_ _1211_ ttA_1.top.backend.wptr_gray\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1706__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ _1142_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2054__S1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3264_ _0227_ net100 ttA_6.counter\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3195_ ttA_1.top.backend.rptr\[3\] _0010_ net38 ttA_1.top.frontend.rptr_gray1\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2131__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2146_ _1083_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _0267_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2434__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2979_ _0893_ _1028_ _1031_ _1007_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2800__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2370__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3288__290 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2189__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3055__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ _1509_ _1343_ _1518_ _1519_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2113__A1 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2902_ _0904_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2833_ _0407_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2764_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1927__A1 ttA_6.counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ _1252_ _1244_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2620__I _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2695_ _0837_ _0838_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1646_ _1165_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1577_ _1129_ _1130_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2352__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3247_ _0210_ net100 ttA_4.active_duty\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3178_ _0158_ net86 ttA_0.data\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2129_ _0350_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3078__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2591__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__S1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2705__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ _1176_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3101_ _0081_ net115 ttA_0.data\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3032_ _1283_ _1059_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3220__CLK net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ ttA_0.data\[2\]\[1\] _0920_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ ttA_0.data\[12\]\[3\] _0873_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2678_ _0735_ _0704_ _0803_ _0822_ _0823_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1629_ _1147_ _1157_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2628__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2100__I1 ttA_0.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2316__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2601_ _0748_ _0739_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2532_ _1223_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2555__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2463_ _0554_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1942__C _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2394_ _0428_ _0572_ _0578_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1530__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3015_ ttA_6.counter\[10\] _1053_ _1346_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout42_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3116__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout110 net117 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xuser_proj_138 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_149 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2085__I0 ttA_0.data\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1963_ ttA_1.top.data\[3\]\[0\] _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1894_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2776__A1 ttA_0.data\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2515_ ttA_0.prog\[5\]\[2\] _0668_ _0670_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2446_ ttA_0.prog\[9\]\[2\] _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3289__CLK clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2377_ ttA_0.prog\[13\]\[1\] _0564_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3008__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2803__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__A1 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2519__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2678__C _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3280_ _0243_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2930__A1 ttA_4.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1733__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2300_ _0496_ _0509_ _0511_ _0507_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2231_ _0448_ _0458_ _0461_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2162_ _0350_ _0409_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_113_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2093_ _1418_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2995_ ttA_6.counter\[4\] _1437_ _1036_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1946_ _1453_ _1468_ _1364_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _1168_ _1078_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1724__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2429_ ttA_0.prog\[10\]\[2\] _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1660__A1 ttA_1.top.backend.wptr_gray\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2912__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2979__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1651__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ _1326_ _1328_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2780_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ _1163_ _1165_ _1166_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ ttA_1.top.frontend.wptr\[2\] ttA_1.top.frontend.wptr\[1\] _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1593_ _1147_ _1129_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2903__A1 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3263_ _0226_ net121 ttA_6.counter\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3194_ ttA_1.top.backend.rptr_b2g.gray\[2\] _0009_ net39 ttA_1.top.frontend.rptr_gray1\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2214_ _1225_ _1226_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2145_ _0381_ _0395_ _0396_ _0390_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2682__A3 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2076_ _0258_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1642__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ ttA_0.data\[11\]\[1\] _1029_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2198__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _1345_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2370__A2 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2122__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2263__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2361__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1624__A1 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ _0977_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2832_ _0927_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2763_ _0476_ _0517_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1714_ _1234_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2901__I _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2694_ _1509_ _0728_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _1152_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1576_ _1105_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3246_ _0209_ net99 ttA_4.active_duty\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout72_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3177_ _0157_ net86 ttA_0.data\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1863__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2128_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2059_ _0291_ _0302_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1615__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2591__A2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2343__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1854__A1 ttA_4.pwm_signal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__B2 ttA_2.io_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__A1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2877__B _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3100_ _0080_ net114 ttA_0.data\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3031_ _0961_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ _0888_ _0919_ _0921_ _0897_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _0857_ _0872_ _0876_ _0877_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2677_ _0389_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1628_ _1160_ _1162_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3462__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1559_ _1099_ _1112_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2089__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3229_ _0192_ net58 ttA_0.prog\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__I _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout122_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _0741_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2531_ _0546_ _0675_ _0680_ _0682_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2462_ _1123_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2393_ ttA_0.prog\[12\]\[2\] _0573_ _0576_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3014_ _1035_ _1054_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout35_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2729_ _0849_ _0864_ _0866_ _0859_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout122 net124 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout100 net101 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_121_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout111 net116 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2482__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_proj_128 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_139 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2085__I1 ttA_0.data\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2537__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ _1252_ ttA_1.top.data\[0\]\[0\] _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1893_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2181__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2514_ _0423_ _0667_ _0671_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1525__I _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2445_ _0616_ _0613_ _0618_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2376_ _0555_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2091__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3233__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2455__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2207__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2066__S0 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ ttA_1.top.data\[2\]\[2\] _0457_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2694__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _1333_ _0345_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2092_ _0313_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2176__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2994_ _1039_ _1040_ _1041_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1945_ _1444_ _1465_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3106__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ net95 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3256__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1724__A3 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ _0603_ _0600_ _0605_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2685__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2359_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2988__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1660__A2 ttA_1.top.frontend.wptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2676__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3129__CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2724__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3279__CLK clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ ttA_2.io_out\[0\] _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _1210_ ttA_1.top.backend.wptr_gray\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1592_ ttA_2.io_out\[6\] _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2903__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3262_ _0225_ net120 ttA_6.counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input7_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2213_ _0448_ _0444_ _0449_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3193_ ttA_1.top.backend.rptr_b2g.gray\[1\] _0008_ net39 ttA_1.top.frontend.rptr_gray1\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2667__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__I _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2144_ ttA_0.data\[1\]\[1\] _0387_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2419__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ _0256_ _0314_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ _0888_ _1028_ _1030_ _1007_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ _1388_ _1446_ _1449_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1859_ ttA_6.counter\[0\] _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2809__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2719__I _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2900_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1624__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__A1 ttA_0.data\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2831_ _0927_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ _0385_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1713_ _1251_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2693_ _0402_ _0748_ _0779_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1644_ _1190_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ ttA_2.io_out\[1\] _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3245_ _0208_ net100 ttA_4.active_duty\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout65_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3176_ _0156_ net88 ttA_0.data\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2127_ _0348_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2058_ _0304_ _0306_ _0308_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2112__I0 ttA_0.data\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1615__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1708__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1551__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2031__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2877__C _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1542__A1 ttA_2.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3030_ _0962_ _1060_ _1061_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2184__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2814_ ttA_0.data\[2\]\[0\] _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2745_ _0681_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2676_ _0756_ _0808_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1781__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _1164_ _1173_ _1175_ _1179_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1558_ ttA_2.io_out\[3\] _1092_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2359__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3228_ _0191_ net57 ttA_0.prog\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3159_ _0139_ net123 ttA_0.io_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2269__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout115_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2461_ ttA_0.prog\[8\]\[1\] _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2392_ _0423_ _0572_ _0577_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _1435_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1967__B _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout28_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2243__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ ttA_0.data\[3\]\[0\] _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2951__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2659_ ttA_0.io_out\[4\] _0342_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout101 net102 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout112 net115 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_129 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_1_1__f_wb_clk_i clknet_0_wb_clk_i clknet_1_1__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2085__I2 ttA_0.data\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1993__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__B _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2170__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _1481_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2462__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1892_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2513_ ttA_0.prog\[5\]\[1\] _0668_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2444_ _0452_ _0614_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2375_ _0549_ _0563_ _0565_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3185__CLK net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1727__B2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1727__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1716__I _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2455__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1966__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1718__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2066__S1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1626__I _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3058__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A1 ttA_0.prog\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2694__A2 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _0359_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2091_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2993_ _1385_ _1037_ _1358_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1944_ _1346_ _1360_ _1388_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2749__A3 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1875_ _1127_ _1076_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1709__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1536__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1724__A4 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _0452_ _0601_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _1370_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2685__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2289_ _0399_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2437__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2988__A3 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2830__I _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3200__CLK net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__B1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2428__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ ttA_1.top.backend.wptr_gray\[3\] ttA_1.top.frontend.wptr\[2\] _1210_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ _1141_ _1143_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3261_ _0224_ net120 ttA_6.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2212_ ttA_1.top.data\[4\]\[2\] _0443_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3192_ ttA_1.top.backend.rptr_b2g.gray\[0\] _0007_ net47 ttA_1.top.frontend.rptr_gray1\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2667__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2143_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2419__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2074_ _0315_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1627__B1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2976_ ttA_0.data\[11\]\[0\] _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1927_ ttA_6.counter\[11\] ttA_6.counter\[10\] ttA_6.counter\[9\] _1450_ _1451_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1858_ ttA_6.counter\[2\] _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1789_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2355__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2658__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2346__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2649__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3246__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2830_ _0927_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2761_ _0860_ _0880_ _0887_ _0886_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1712_ _1250_ ttA_1.top.backend.rptr_b2g.gray\[0\] _1244_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2692_ _0402_ _0748_ _0757_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1643_ _1097_ _1114_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3244_ _0207_ net94 ttA_4.active_duty\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3175_ _0155_ net104 ttA_0.data\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1863__A3 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2126_ _0349_ _0364_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_fanout58_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2057_ _0297_ _0309_ _0255_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2112__I1 ttA_0.data\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2959_ _1368_ _1015_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2328__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3269__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2983__C _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1599__C _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__A1 ttA_0.data\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1542__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ _0918_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__S0 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2744_ ttA_0.data\[12\]\[2\] _0873_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2675_ _0767_ _0815_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1626_ _1159_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1557_ _1107_ _1110_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2730__A1 ttA_0.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3227_ _0190_ net52 ttA_0.prog\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3158_ _0138_ net118 ttA_0.io_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2109_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_0__f_wb_clk_i clknet_0_wb_clk_i clknet_1_0__leaf_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3089_ _0069_ net109 ttA_0.data\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2564__A4 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3091__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2960__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _0625_ _0628_ _0630_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2391_ ttA_0.prog\[12\]\[1\] _0573_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3012_ _0960_ _1052_ _1053_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1967__C _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2779__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ _0863_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2951__B2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2951__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ _0734_ _0361_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout102 net126 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1609_ _1089_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2589_ _1508_ _0409_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout113 net114 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_102_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2833__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2942__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1960_ ttA_1.top.data\[1\]\[0\] _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2512_ _0633_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2933__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2443_ _0575_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2374_ ttA_0.prog\[13\]\[0\] _0564_ _0557_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout40_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1978__B _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2915__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__I ttA_0.io_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1798__B _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2473__I ttA_0.prog\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2992_ _1438_ _1037_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1943_ _1358_ _1385_ _1447_ _1448_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1874_ _1370_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1817__I _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2906__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2382__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2426_ _0575_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3152__CLK net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout88_I net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0551_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2288_ _0501_ _0498_ _0502_ _0495_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2070__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1590_ _1144_ _1143_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2364__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3260_ _0223_ net119 ttA_6.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _1160_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3191_ ttA_1.top.frontend.rptr_gray1\[3\] _0006_ net38 ttA_1.top.frontend.rptr_gray2\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_121_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1875__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2142_ _0392_ _0382_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2073_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1975__C _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2975_ _1027_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xuser_proj_280 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1926_ ttA_6.counter\[8\] _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1857_ _1334_ _1343_ _1384_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ beepboop.inst.counter\[3\] beepboop.inst.counter\[2\] _1275_ _1317_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2409_ _0588_ _0584_ _0590_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2291__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3198__CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1857__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2751__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2760_ ttA_0.data\[15\]\[3\] _0881_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1711_ _1233_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2691_ _0737_ _0829_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1642_ _1190_ _1184_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1573_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3243_ _0206_ net97 ttA_4.active_duty\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ _0154_ net104 ttA_0.data\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1830__I ttA_6.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2125_ _0375_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2056_ ttA_0.prog\[4\]\[1\] ttA_0.prog\[5\]\[1\] ttA_0.prog\[6\]\[1\] ttA_0.prog\[7\]\[1\]
+ _0298_ _0299_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2112__I2 ttA_0.data\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2958_ _1402_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2576__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1909_ _1432_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2889_ ttA_0.prog\[1\]\[1\] _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2836__I ttA_4.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2057__B _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2264__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3213__CLK net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2481__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2812_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2558__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2102__S1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2743_ _0855_ _0872_ _0875_ _0869_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2674_ _0817_ _0818_ _0819_ _0754_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1625_ _1176_ _1178_ _1123_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1556_ ttA_2.io_out\[2\] _1109_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout70_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3226_ _0189_ net57 ttA_0.prog\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3157_ _0137_ net109 ttA_0.io_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2494__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2108_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3088_ _0068_ net112 ttA_0.data\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2246__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ ttA_0.io_out\[2\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1735__I _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3236__CLK net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2515__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2390_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3011_ _1441_ _1051_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2476__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3109__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__S0 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2726_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2951__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _0796_ _0799_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1608_ ttA_2.io_out\[6\] _1094_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2588_ _0409_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout103 net105 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout125 net126 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1539_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3209_ ttA_1.top.backend.wptr_gray\[1\] _0020_ net28 ttA_1.top.backend.wptr_gray1\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2011__S0 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2219__A1 ttA_1.top.data\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__S0 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2630__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1890_ ttA_0.io_out\[2\] _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2069__S0 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout120_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2511_ _0534_ _0667_ _0669_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2933__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2442_ ttA_0.prog\[9\]\[1\] _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2697__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2373_ _0562_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2934__I _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2709_ _0851_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2860__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2915__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1923__I _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2679__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ _0959_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1942_ _1436_ _1459_ _1464_ _1443_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ _1366_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2906__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1590__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2425_ ttA_0.prog\[10\]\[1\] _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2287_ ttA_0.data\[8\]\[1\] _0499_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A2 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1581__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2839__I ttA_4.active_duty\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1636__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0446_ _0444_ _0447_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3190_ ttA_1.top.frontend.rptr_gray1\[2\] _0005_ net38 ttA_1.top.frontend.rptr_gray2\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_121_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2141_ _1153_ _0383_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2072_ _0317_ _0320_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2974_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1925_ _1447_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xuser_proj_270 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_281 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1856_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1787_ _1284_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2408_ _0452_ _0586_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2339_ _1419_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I io_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1618__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2815__A1 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2043__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1554__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3142__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1710_ _1249_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2690_ _0830_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1641_ _1193_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ _1091_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2479__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3242_ _0205_ net85 ttA_0.data\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3173_ _0153_ net106 ttA_0.data\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2124_ _0376_ _0315_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2055_ _1417_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2957_ ttA_0.lastdata3 _0700_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2025__A2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1908_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2888_ _0964_ _0966_ _0969_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1839_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2389__I _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3165__CLK net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A3 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2762__I _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2811_ _0348_ _0517_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ ttA_0.data\[12\]\[1\] _0873_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _0778_ _0749_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1624_ _1141_ _1166_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ ttA_2.io_out\[2\] _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3225_ _0188_ net57 ttA_0.prog\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1841__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _0136_ net75 ttA_1.top.data\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout63_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__A2 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2107_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3087_ _0067_ net109 ttA_0.data\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2038_ _0286_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2246__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1757__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__A1 ttA_1.top.data\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1996__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2757__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3010_ _1441_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__S1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1836__I _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2400__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2725_ _0348_ _0485_ _0486_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2656_ _0796_ _0799_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1607_ _1096_ _1118_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2587_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2164__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout104 net107 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout126 net127 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_141_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1538_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout115 net116 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1571__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3208_ ttA_1.top.backend.wptr_gray\[0\] _0019_ net29 ttA_1.top.backend.wptr_gray1\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2011__S1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3139_ _0119_ net54 ttA_0.prog\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1978__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3203__CLK net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2078__S1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1745__A4 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__A1 _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1902__B2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2069__S1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2394__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout113_I net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2510_ ttA_0.prog\[5\]\[0\] _0668_ _0662_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2441_ _0610_ _0613_ _0615_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2697__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2372_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2449__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3226__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2950__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2621__A2 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2639_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2688__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3021__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2679__A2 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3249__CLK net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2300__A1 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2990_ _1035_ _1038_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1941_ _1441_ _1436_ _1389_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1872_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2367__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A2 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _0597_ _0600_ _0602_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2355_ _0550_ _0539_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2286_ _0394_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2855__I ttA_0.prog\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2523__C _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3071__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2140_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _0287_ _0321_ _0323_ _0256_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2765__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0485_ _0486_ _0476_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_proj_260 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1924_ ttA_6.counter\[4\] _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_proj_271 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xuser_proj_282 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1855_ _1356_ _1365_ _1367_ _1379_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_135_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1786_ beepboop.inst.counter\[10\] _1306_ beepboop.inst.counter\[8\] _1315_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1844__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2407_ _0575_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2338_ _0256_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2269_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2624__B _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2579__B2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3158__D _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2585__I _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2114__S0 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2990__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1640_ _1192_ _1144_ _1085_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1571_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2742__A1 ttA_0.data\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3241_ _0204_ net82 ttA_0.data\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3172_ _0152_ net106 ttA_0.data\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ _1396_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2054_ ttA_0.prog\[0\]\[1\] ttA_0.prog\[1\]\[1\] ttA_0.prog\[2\]\[1\] ttA_0.prog\[3\]\[1\]
+ _0293_ _0294_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2956_ _1376_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1907_ ttA_0.io_out\[3\] _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2887_ _0647_ _0967_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1838_ net9 _1339_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2981__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1769_ _1289_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1749__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2972__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1659__I ttA_1.top.frontend.wptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2810_ _0917_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2741_ _0849_ _0872_ _0874_ _0869_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2963__A1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _0735_ _0816_ _0736_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2711__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ ttA_2.io_out\[3\] _1168_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1554_ net6 _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3224_ _0187_ clknet_1_0__leaf_wb_clk_i beepboop.inst.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends


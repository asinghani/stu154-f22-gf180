// This is the unpowered netlist.
module user_proj (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire net295;
 wire net294;
 wire net293;
 wire net292;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire net291;
 wire net290;
 wire net289;
 wire net288;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire \beepboop.inst.counter[0] ;
 wire \beepboop.inst.counter[10] ;
 wire \beepboop.inst.counter[11] ;
 wire \beepboop.inst.counter[12] ;
 wire \beepboop.inst.counter[13] ;
 wire \beepboop.inst.counter[14] ;
 wire \beepboop.inst.counter[15] ;
 wire \beepboop.inst.counter[1] ;
 wire \beepboop.inst.counter[2] ;
 wire \beepboop.inst.counter[3] ;
 wire \beepboop.inst.counter[4] ;
 wire \beepboop.inst.counter[5] ;
 wire \beepboop.inst.counter[6] ;
 wire \beepboop.inst.counter[7] ;
 wire \beepboop.inst.counter[8] ;
 wire \beepboop.inst.counter[9] ;
 wire net129;
 wire net296;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net297;
 wire net146;
 wire net130;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net131;
 wire clknet_0_wb_clk_i;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net164;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net165;
 wire net184;
 wire net185;
 wire net166;
 wire net186;
 wire net187;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net192;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net193;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net194;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net195;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net196;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire \ttA_0.data[0][0] ;
 wire \ttA_0.data[0][1] ;
 wire \ttA_0.data[0][2] ;
 wire \ttA_0.data[0][3] ;
 wire \ttA_0.data[10][0] ;
 wire \ttA_0.data[10][1] ;
 wire \ttA_0.data[10][2] ;
 wire \ttA_0.data[10][3] ;
 wire \ttA_0.data[11][0] ;
 wire \ttA_0.data[11][1] ;
 wire \ttA_0.data[11][2] ;
 wire \ttA_0.data[11][3] ;
 wire \ttA_0.data[12][0] ;
 wire \ttA_0.data[12][1] ;
 wire \ttA_0.data[12][2] ;
 wire \ttA_0.data[12][3] ;
 wire \ttA_0.data[13][0] ;
 wire \ttA_0.data[13][1] ;
 wire \ttA_0.data[13][2] ;
 wire \ttA_0.data[13][3] ;
 wire \ttA_0.data[14][0] ;
 wire \ttA_0.data[14][1] ;
 wire \ttA_0.data[14][2] ;
 wire \ttA_0.data[14][3] ;
 wire \ttA_0.data[15][0] ;
 wire \ttA_0.data[15][1] ;
 wire \ttA_0.data[15][2] ;
 wire \ttA_0.data[15][3] ;
 wire \ttA_0.data[1][0] ;
 wire \ttA_0.data[1][1] ;
 wire \ttA_0.data[1][2] ;
 wire \ttA_0.data[1][3] ;
 wire \ttA_0.data[2][0] ;
 wire \ttA_0.data[2][1] ;
 wire \ttA_0.data[2][2] ;
 wire \ttA_0.data[2][3] ;
 wire \ttA_0.data[3][0] ;
 wire \ttA_0.data[3][1] ;
 wire \ttA_0.data[3][2] ;
 wire \ttA_0.data[3][3] ;
 wire \ttA_0.data[4][0] ;
 wire \ttA_0.data[4][1] ;
 wire \ttA_0.data[4][2] ;
 wire \ttA_0.data[4][3] ;
 wire \ttA_0.data[5][0] ;
 wire \ttA_0.data[5][1] ;
 wire \ttA_0.data[5][2] ;
 wire \ttA_0.data[5][3] ;
 wire \ttA_0.data[6][0] ;
 wire \ttA_0.data[6][1] ;
 wire \ttA_0.data[6][2] ;
 wire \ttA_0.data[6][3] ;
 wire \ttA_0.data[7][0] ;
 wire \ttA_0.data[7][1] ;
 wire \ttA_0.data[7][2] ;
 wire \ttA_0.data[7][3] ;
 wire \ttA_0.data[8][0] ;
 wire \ttA_0.data[8][1] ;
 wire \ttA_0.data[8][2] ;
 wire \ttA_0.data[8][3] ;
 wire \ttA_0.data[9][0] ;
 wire \ttA_0.data[9][1] ;
 wire \ttA_0.data[9][2] ;
 wire \ttA_0.data[9][3] ;
 wire \ttA_0.io_out[0] ;
 wire \ttA_0.io_out[1] ;
 wire \ttA_0.io_out[2] ;
 wire \ttA_0.io_out[3] ;
 wire \ttA_0.io_out[4] ;
 wire \ttA_0.io_out[5] ;
 wire \ttA_0.io_out[6] ;
 wire \ttA_0.io_out[7] ;
 wire \ttA_0.lastdata3 ;
 wire \ttA_0.prog[0][0] ;
 wire \ttA_0.prog[0][1] ;
 wire \ttA_0.prog[0][2] ;
 wire \ttA_0.prog[0][3] ;
 wire \ttA_0.prog[10][0] ;
 wire \ttA_0.prog[10][1] ;
 wire \ttA_0.prog[10][2] ;
 wire \ttA_0.prog[10][3] ;
 wire \ttA_0.prog[11][0] ;
 wire \ttA_0.prog[11][1] ;
 wire \ttA_0.prog[11][2] ;
 wire \ttA_0.prog[11][3] ;
 wire \ttA_0.prog[12][0] ;
 wire \ttA_0.prog[12][1] ;
 wire \ttA_0.prog[12][2] ;
 wire \ttA_0.prog[12][3] ;
 wire \ttA_0.prog[13][0] ;
 wire \ttA_0.prog[13][1] ;
 wire \ttA_0.prog[13][2] ;
 wire \ttA_0.prog[13][3] ;
 wire \ttA_0.prog[14][0] ;
 wire \ttA_0.prog[14][1] ;
 wire \ttA_0.prog[14][2] ;
 wire \ttA_0.prog[14][3] ;
 wire \ttA_0.prog[15][0] ;
 wire \ttA_0.prog[15][1] ;
 wire \ttA_0.prog[15][2] ;
 wire \ttA_0.prog[15][3] ;
 wire \ttA_0.prog[1][0] ;
 wire \ttA_0.prog[1][1] ;
 wire \ttA_0.prog[1][2] ;
 wire \ttA_0.prog[1][3] ;
 wire \ttA_0.prog[2][0] ;
 wire \ttA_0.prog[2][1] ;
 wire \ttA_0.prog[2][2] ;
 wire \ttA_0.prog[2][3] ;
 wire \ttA_0.prog[3][0] ;
 wire \ttA_0.prog[3][1] ;
 wire \ttA_0.prog[3][2] ;
 wire \ttA_0.prog[3][3] ;
 wire \ttA_0.prog[4][0] ;
 wire \ttA_0.prog[4][1] ;
 wire \ttA_0.prog[4][2] ;
 wire \ttA_0.prog[4][3] ;
 wire \ttA_0.prog[5][0] ;
 wire \ttA_0.prog[5][1] ;
 wire \ttA_0.prog[5][2] ;
 wire \ttA_0.prog[5][3] ;
 wire \ttA_0.prog[6][0] ;
 wire \ttA_0.prog[6][1] ;
 wire \ttA_0.prog[6][2] ;
 wire \ttA_0.prog[6][3] ;
 wire \ttA_0.prog[7][0] ;
 wire \ttA_0.prog[7][1] ;
 wire \ttA_0.prog[7][2] ;
 wire \ttA_0.prog[7][3] ;
 wire \ttA_0.prog[8][0] ;
 wire \ttA_0.prog[8][1] ;
 wire \ttA_0.prog[8][2] ;
 wire \ttA_0.prog[8][3] ;
 wire \ttA_0.prog[9][0] ;
 wire \ttA_0.prog[9][1] ;
 wire \ttA_0.prog[9][2] ;
 wire \ttA_0.prog[9][3] ;
 wire \ttA_1.top.backend.rptr[0] ;
 wire \ttA_1.top.backend.rptr[1] ;
 wire \ttA_1.top.backend.rptr[2] ;
 wire \ttA_1.top.backend.rptr[3] ;
 wire \ttA_1.top.backend.rptr_b2g.gray[0] ;
 wire \ttA_1.top.backend.rptr_b2g.gray[1] ;
 wire \ttA_1.top.backend.rptr_b2g.gray[2] ;
 wire \ttA_1.top.backend.wptr_gray1[0] ;
 wire \ttA_1.top.backend.wptr_gray1[1] ;
 wire \ttA_1.top.backend.wptr_gray1[2] ;
 wire \ttA_1.top.backend.wptr_gray1[3] ;
 wire \ttA_1.top.backend.wptr_gray2[0] ;
 wire \ttA_1.top.backend.wptr_gray2[1] ;
 wire \ttA_1.top.backend.wptr_gray2[2] ;
 wire \ttA_1.top.backend.wptr_gray2[3] ;
 wire \ttA_1.top.backend.wptr_gray[0] ;
 wire \ttA_1.top.backend.wptr_gray[1] ;
 wire \ttA_1.top.backend.wptr_gray[2] ;
 wire \ttA_1.top.backend.wptr_gray[3] ;
 wire \ttA_1.top.data[0][0] ;
 wire \ttA_1.top.data[0][1] ;
 wire \ttA_1.top.data[0][2] ;
 wire \ttA_1.top.data[1][0] ;
 wire \ttA_1.top.data[1][1] ;
 wire \ttA_1.top.data[1][2] ;
 wire \ttA_1.top.data[2][0] ;
 wire \ttA_1.top.data[2][1] ;
 wire \ttA_1.top.data[2][2] ;
 wire \ttA_1.top.data[3][0] ;
 wire \ttA_1.top.data[3][1] ;
 wire \ttA_1.top.data[3][2] ;
 wire \ttA_1.top.data[4][0] ;
 wire \ttA_1.top.data[4][1] ;
 wire \ttA_1.top.data[4][2] ;
 wire \ttA_1.top.data[5][0] ;
 wire \ttA_1.top.data[5][1] ;
 wire \ttA_1.top.data[5][2] ;
 wire \ttA_1.top.data[6][0] ;
 wire \ttA_1.top.data[6][1] ;
 wire \ttA_1.top.data[6][2] ;
 wire \ttA_1.top.data[7][0] ;
 wire \ttA_1.top.data[7][1] ;
 wire \ttA_1.top.data[7][2] ;
 wire \ttA_1.top.frontend.rptr_gray1[0] ;
 wire \ttA_1.top.frontend.rptr_gray1[1] ;
 wire \ttA_1.top.frontend.rptr_gray1[2] ;
 wire \ttA_1.top.frontend.rptr_gray1[3] ;
 wire \ttA_1.top.frontend.rptr_gray2[0] ;
 wire \ttA_1.top.frontend.rptr_gray2[1] ;
 wire \ttA_1.top.frontend.rptr_gray2[2] ;
 wire \ttA_1.top.frontend.rptr_gray2[3] ;
 wire \ttA_1.top.frontend.wptr[0] ;
 wire \ttA_1.top.frontend.wptr[1] ;
 wire \ttA_1.top.frontend.wptr[2] ;
 wire \ttA_2.io_out[0] ;
 wire \ttA_2.io_out[1] ;
 wire \ttA_2.io_out[2] ;
 wire \ttA_2.io_out[3] ;
 wire \ttA_2.io_out[4] ;
 wire \ttA_2.io_out[5] ;
 wire \ttA_2.io_out[6] ;
 wire \ttA_2.io_out[7] ;
 wire \ttA_2.state ;
 wire \ttA_4.active_duty[0] ;
 wire \ttA_4.active_duty[1] ;
 wire \ttA_4.active_duty[2] ;
 wire \ttA_4.active_duty[3] ;
 wire \ttA_4.active_duty[4] ;
 wire \ttA_4.active_duty[5] ;
 wire \ttA_4.counter[0] ;
 wire \ttA_4.counter[1] ;
 wire \ttA_4.counter[2] ;
 wire \ttA_4.counter[3] ;
 wire \ttA_4.counter[4] ;
 wire \ttA_4.counter[5] ;
 wire \ttA_4.pwm_signal ;
 wire \ttA_6.counter[0] ;
 wire \ttA_6.counter[10] ;
 wire \ttA_6.counter[11] ;
 wire \ttA_6.counter[12] ;
 wire \ttA_6.counter[13] ;
 wire \ttA_6.counter[14] ;
 wire \ttA_6.counter[15] ;
 wire \ttA_6.counter[1] ;
 wire \ttA_6.counter[2] ;
 wire \ttA_6.counter[3] ;
 wire \ttA_6.counter[4] ;
 wire \ttA_6.counter[5] ;
 wire \ttA_6.counter[6] ;
 wire \ttA_6.counter[7] ;
 wire \ttA_6.counter[8] ;
 wire \ttA_6.counter[9] ;
 wire net255;
 wire net256;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net257;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net258;
 wire net286;
 wire net287;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1521_ (.I(net3),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1522_ (.I(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1523_ (.I(_1077_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1524_ (.A1(_1078_),
    .A2(\ttA_2.state ),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1525_ (.I(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1526_ (.I(net8),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1527_ (.I(net7),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1528_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1529_ (.A1(_1081_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1530_ (.A1(_1080_),
    .A2(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1531_ (.I(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1532_ (.I(_1081_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1533_ (.I(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1534_ (.I(net6),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1535_ (.I(net5),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1536_ (.I(net4),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1537_ (.A1(_1089_),
    .A2(_1090_),
    .A3(_1091_),
    .B1(_1083_),
    .B2(net8),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1538_ (.I(_1092_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1539_ (.I(_1093_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1540_ (.A1(\ttA_2.io_out[6] ),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1541_ (.A1(\ttA_2.io_out[5] ),
    .A2(_1093_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1542_ (.A1(\ttA_2.io_out[4] ),
    .A2(_1092_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1543_ (.I(\ttA_2.io_out[3] ),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1544_ (.A1(_1098_),
    .A2(_1092_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1545_ (.I(\ttA_2.io_out[1] ),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1546_ (.A1(net8),
    .A2(_1082_),
    .B(net4),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1547_ (.A1(_1090_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1548_ (.A1(_1090_),
    .A2(_1101_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1549_ (.I(_1091_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1550_ (.A1(_1104_),
    .A2(\ttA_2.io_out[0] ),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1551_ (.A1(net5),
    .A2(_1100_),
    .A3(_1101_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1552_ (.A1(_1100_),
    .A2(_1102_),
    .A3(_1103_),
    .B1(_1105_),
    .B2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1553_ (.A1(net8),
    .A2(_1083_),
    .B1(net5),
    .B2(net4),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1554_ (.A1(net6),
    .A2(_1108_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1555_ (.A1(\ttA_2.io_out[2] ),
    .A2(_1109_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1556_ (.A1(\ttA_2.io_out[2] ),
    .A2(_1109_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1557_ (.A1(_1107_),
    .A2(_1110_),
    .B(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1558_ (.A1(\ttA_2.io_out[3] ),
    .A2(_1092_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1559_ (.A1(_1099_),
    .A2(_1112_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1560_ (.A1(\ttA_2.io_out[5] ),
    .A2(_1093_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(\ttA_2.io_out[4] ),
    .A2(_1093_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1562_ (.I(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1563_ (.A1(_1097_),
    .A2(_1114_),
    .B(_1115_),
    .C(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1564_ (.A1(\ttA_2.io_out[6] ),
    .A2(_1094_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1565_ (.A1(_1095_),
    .A2(_1096_),
    .A3(_1118_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1566_ (.A1(\ttA_2.io_out[7] ),
    .A2(_1094_),
    .A3(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1567_ (.I(_1087_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1568_ (.I(_1089_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1569_ (.I(_1090_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1570_ (.I(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1571_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1572_ (.I(_1091_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1573_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1574_ (.I(_1128_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1575_ (.I(\ttA_2.io_out[1] ),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1576_ (.I(_1105_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1577_ (.A1(_1129_),
    .A2(_1130_),
    .B(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1578_ (.I(_1125_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1579_ (.I(\ttA_2.io_out[2] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1580_ (.A1(_1128_),
    .A2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1581_ (.A1(_1098_),
    .A2(_1128_),
    .B(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1582_ (.A1(_1133_),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1583_ (.A1(_1126_),
    .A2(_1132_),
    .B(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1584_ (.A1(_1123_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1585_ (.I(_1133_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1586_ (.I(\ttA_2.io_out[4] ),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1587_ (.I(_1104_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1588_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1589_ (.I(\ttA_2.io_out[5] ),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1590_ (.A1(_1144_),
    .A2(_1143_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1591_ (.A1(_1141_),
    .A2(_1143_),
    .B(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1592_ (.I(\ttA_2.io_out[6] ),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(_1147_),
    .A2(_1129_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1594_ (.I(_1142_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1595_ (.A1(\ttA_2.io_out[7] ),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1596_ (.A1(_1126_),
    .A2(_1148_),
    .A3(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1597_ (.I(_1089_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1598_ (.I(_1152_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1599_ (.A1(_1140_),
    .A2(_1146_),
    .B(_1151_),
    .C(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1600_ (.A1(_1122_),
    .A2(_1139_),
    .A3(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1601_ (.A1(_1088_),
    .A2(_1121_),
    .B(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1602_ (.I(_1085_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1603_ (.A1(\ttA_2.io_out[7] ),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1604_ (.A1(_1086_),
    .A2(_1156_),
    .B(_1158_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1605_ (.I(_1081_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1606_ (.I(_1159_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1607_ (.A1(_1096_),
    .A2(_1118_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1608_ (.A1(\ttA_2.io_out[6] ),
    .A2(_1094_),
    .A3(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1609_ (.I(_1089_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1610_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1611_ (.I(_1124_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1612_ (.I(_1128_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1613_ (.I(_1134_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1614_ (.I(_1127_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1615_ (.A1(_1168_),
    .A2(_1130_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1616_ (.A1(_1166_),
    .A2(_1167_),
    .B(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1617_ (.A1(_1143_),
    .A2(\ttA_2.io_out[0] ),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1618_ (.A1(_1124_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1619_ (.A1(_1165_),
    .A2(_1170_),
    .B(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1620_ (.A1(_1147_),
    .A2(_1129_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1621_ (.A1(_1144_),
    .A2(_1149_),
    .B(_1174_),
    .C(_1126_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1622_ (.I(_1124_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(\ttA_2.io_out[3] ),
    .A2(_1168_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1624_ (.A1(_1141_),
    .A2(_1166_),
    .B(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1625_ (.A1(_1176_),
    .A2(_1178_),
    .B(_1123_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1626_ (.I(_1159_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1627_ (.A1(_1164_),
    .A2(_1173_),
    .B1(_1175_),
    .B2(_1179_),
    .C(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1628_ (.A1(_1160_),
    .A2(_1162_),
    .B(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1629_ (.A1(_1147_),
    .A2(_1157_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(_1086_),
    .A2(_1182_),
    .B(_1183_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1631_ (.A1(_1097_),
    .A2(_1114_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1632_ (.A1(_1117_),
    .A2(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1633_ (.A1(_1115_),
    .A2(_1096_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1634_ (.A1(_1185_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1635_ (.I0(_1136_),
    .I1(_1146_),
    .S(_1133_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1636_ (.A1(_1165_),
    .A2(_1132_),
    .B(_1163_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1637_ (.I(_1081_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1638_ (.A1(_1164_),
    .A2(_1188_),
    .B(_1189_),
    .C(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1639_ (.A1(_1122_),
    .A2(_1187_),
    .B(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1640_ (.I0(_1192_),
    .I1(_1144_),
    .S(_1085_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1641_ (.I(_1193_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1642_ (.A1(_1190_),
    .A2(_1184_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1643_ (.A1(_1097_),
    .A2(_1114_),
    .B(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1644_ (.I(_1190_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1645_ (.I(_1152_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1646_ (.I(_1165_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1647_ (.A1(_1140_),
    .A2(_1170_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1648_ (.A1(_1176_),
    .A2(_1178_),
    .B(_1153_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1649_ (.A1(_1197_),
    .A2(_1198_),
    .A3(_1171_),
    .B1(_1199_),
    .B2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1650_ (.A1(_1196_),
    .A2(_1201_),
    .B(_1157_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1651_ (.A1(_1141_),
    .A2(_1086_),
    .B1(_1195_),
    .B2(_1202_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1652_ (.A1(_1099_),
    .A2(_1112_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1653_ (.A1(_1160_),
    .A2(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1654_ (.I(_1163_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1655_ (.A1(_1180_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1656_ (.A1(_1138_),
    .A2(_1206_),
    .B(_1157_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1657_ (.A1(_1098_),
    .A2(_1086_),
    .B1(_1204_),
    .B2(_1207_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1658_ (.I(\ttA_1.top.frontend.wptr[2] ),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1659_ (.I(\ttA_1.top.frontend.wptr[1] ),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1660_ (.A1(\ttA_1.top.backend.wptr_gray[3] ),
    .A2(\ttA_1.top.frontend.wptr[2] ),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1661_ (.I(_1210_),
    .Z(\ttA_1.top.backend.wptr_gray[2] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1662_ (.A1(\ttA_1.top.frontend.wptr[2] ),
    .A2(\ttA_1.top.frontend.wptr[1] ),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1663_ (.I(_1211_),
    .Z(\ttA_1.top.backend.wptr_gray[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1664_ (.I(\ttA_1.top.frontend.rptr_gray2[1] ),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1665_ (.A1(\ttA_1.top.frontend.rptr_gray2[2] ),
    .A2(\ttA_1.top.backend.wptr_gray[2] ),
    .B1(\ttA_1.top.backend.wptr_gray[1] ),
    .B2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1666_ (.A1(\ttA_1.top.frontend.rptr_gray2[2] ),
    .A2(\ttA_1.top.backend.wptr_gray[2] ),
    .B(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1667_ (.A1(\ttA_1.top.frontend.wptr[1] ),
    .A2(\ttA_1.top.frontend.wptr[0] ),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1668_ (.I(_1215_),
    .Z(\ttA_1.top.backend.wptr_gray[0] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1669_ (.A1(\ttA_1.top.frontend.rptr_gray2[0] ),
    .A2(\ttA_1.top.backend.wptr_gray[0] ),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1670_ (.A1(\ttA_1.top.backend.wptr_gray[3] ),
    .A2(\ttA_1.top.frontend.rptr_gray2[3] ),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1671_ (.A1(_1212_),
    .A2(\ttA_1.top.backend.wptr_gray[1] ),
    .B(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1672_ (.A1(_1214_),
    .A2(_1216_),
    .A3(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1673_ (.I(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1674_ (.A1(_1142_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1675_ (.A1(\ttA_1.top.frontend.wptr[0] ),
    .A2(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1676_ (.A1(_1208_),
    .A2(_1209_),
    .A3(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1677_ (.A1(\ttA_1.top.backend.wptr_gray[3] ),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1678_ (.I(_1224_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1679_ (.I(\ttA_1.top.frontend.wptr[2] ),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1680_ (.A1(_1209_),
    .A2(_1222_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1681_ (.A1(_1225_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1682_ (.I(_1227_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1683_ (.I(\ttA_1.top.frontend.wptr[1] ),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1684_ (.A1(\ttA_1.top.backend.wptr_gray[0] ),
    .A2(_1221_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1685_ (.A1(_1228_),
    .A2(_1221_),
    .B(_1229_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1686_ (.A1(\ttA_1.top.frontend.wptr[0] ),
    .A2(_1221_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1687_ (.I(_1230_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1688_ (.I(\ttA_1.top.backend.rptr[2] ),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1689_ (.A1(\ttA_1.top.backend.rptr[3] ),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1690_ (.I(\ttA_1.top.backend.rptr[1] ),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1691_ (.I(\ttA_1.top.backend.rptr[0] ),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1692_ (.I(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1693_ (.A1(\ttA_1.top.backend.rptr[2] ),
    .A2(\ttA_1.top.backend.rptr[1] ),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1694_ (.I(_1236_),
    .Z(\ttA_1.top.backend.rptr_b2g.gray[1] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1695_ (.A1(\ttA_1.top.backend.wptr_gray2[1] ),
    .A2(\ttA_1.top.backend.rptr_b2g.gray[1] ),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1696_ (.A1(\ttA_1.top.backend.rptr[1] ),
    .A2(\ttA_1.top.backend.rptr[0] ),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1697_ (.I(_1238_),
    .Z(\ttA_1.top.backend.rptr_b2g.gray[0] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1698_ (.A1(\ttA_1.top.backend.wptr_gray2[0] ),
    .A2(\ttA_1.top.backend.rptr_b2g.gray[0] ),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1699_ (.A1(\ttA_1.top.backend.wptr_gray2[2] ),
    .A2(_1232_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1700_ (.A1(\ttA_1.top.backend.rptr[3] ),
    .A2(\ttA_1.top.backend.wptr_gray2[3] ),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1701_ (.A1(\ttA_1.top.backend.wptr_gray2[2] ),
    .A2(_1232_),
    .B(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1702_ (.A1(_1237_),
    .A2(_1239_),
    .A3(_1240_),
    .A4(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1703_ (.A1(_1125_),
    .A2(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1704_ (.A1(_1233_),
    .A2(_1235_),
    .A3(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1705_ (.A1(\ttA_1.top.backend.rptr[2] ),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1706_ (.A1(_1232_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1707_ (.I(_1247_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1708_ (.I(_1231_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1709_ (.A1(_1248_),
    .A2(_1245_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1710_ (.I(_1249_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1711_ (.I(_1233_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1712_ (.I0(_1250_),
    .I1(\ttA_1.top.backend.rptr_b2g.gray[0] ),
    .S(_1244_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1713_ (.I(_1251_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1714_ (.I(_1234_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1715_ (.A1(_1252_),
    .A2(_1244_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1716_ (.I(_1253_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1717_ (.A1(_1153_),
    .A2(_1134_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1718_ (.A1(_1084_),
    .A2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1719_ (.A1(_1087_),
    .A2(net7),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1720_ (.A1(_1167_),
    .A2(_1109_),
    .A3(_1107_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1721_ (.A1(_1164_),
    .A2(_1173_),
    .A3(_1256_),
    .B1(_1257_),
    .B2(_1122_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1722_ (.A1(_1255_),
    .A2(_1258_),
    .B(_1080_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1723_ (.A1(_1167_),
    .A2(_1080_),
    .B(_1259_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1724_ (.A1(_1164_),
    .A2(_1198_),
    .A3(_1132_),
    .A4(_1256_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1725_ (.A1(_1131_),
    .A2(_1106_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1726_ (.A1(_1133_),
    .A2(_1130_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1727_ (.A1(_1190_),
    .A2(_1261_),
    .B1(_1262_),
    .B2(_1084_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1728_ (.A1(_1079_),
    .A2(_1260_),
    .A3(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1729_ (.A1(_1100_),
    .A2(_1079_),
    .B(_1264_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1730_ (.I(\ttA_2.io_out[0] ),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1731_ (.A1(_1163_),
    .A2(_1165_),
    .A3(_1166_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1732_ (.A1(_1079_),
    .A2(_1131_),
    .B(_1171_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1733_ (.A1(_1266_),
    .A2(_1256_),
    .B(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1734_ (.A1(_1265_),
    .A2(_1080_),
    .B(_1268_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1735_ (.I(_1232_),
    .ZN(\ttA_1.top.backend.rptr_b2g.gray[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1736_ (.A1(\beepboop.inst.counter[10] ),
    .A2(\beepboop.inst.counter[9] ),
    .A3(\beepboop.inst.counter[8] ),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1737_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1738_ (.A1(\beepboop.inst.counter[15] ),
    .A2(\beepboop.inst.counter[14] ),
    .A3(\beepboop.inst.counter[13] ),
    .A4(\beepboop.inst.counter[12] ),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1739_ (.A1(\beepboop.inst.counter[11] ),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1740_ (.I(\beepboop.inst.counter[2] ),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1741_ (.I(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1742_ (.I(\beepboop.inst.counter[5] ),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1743_ (.I(\beepboop.inst.counter[3] ),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1744_ (.A1(\beepboop.inst.counter[7] ),
    .A2(\beepboop.inst.counter[6] ),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1745_ (.A1(_1275_),
    .A2(\beepboop.inst.counter[4] ),
    .A3(_1276_),
    .A4(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1746_ (.A1(\beepboop.inst.counter[1] ),
    .A2(\beepboop.inst.counter[0] ),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1747_ (.A1(_1274_),
    .A2(_1278_),
    .A3(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1748_ (.A1(_1270_),
    .A2(_1272_),
    .A3(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1749_ (.I(_1271_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1750_ (.A1(\beepboop.inst.counter[4] ),
    .A2(\beepboop.inst.counter[3] ),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1751_ (.I(\beepboop.inst.counter[7] ),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1752_ (.A1(\beepboop.inst.counter[6] ),
    .A2(_1275_),
    .A3(_1283_),
    .B(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1753_ (.A1(_1269_),
    .A2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1754_ (.A1(\beepboop.inst.counter[11] ),
    .A2(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1755_ (.A1(_1282_),
    .A2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1756_ (.I(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1757_ (.A1(_1281_),
    .A2(_1289_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1758_ (.I(_1275_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1759_ (.I(_1290_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1760_ (.I(\beepboop.inst.counter[4] ),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1761_ (.I(_1292_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1762_ (.A1(_1291_),
    .A2(_1293_),
    .A3(_1276_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1763_ (.I(_1284_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1764_ (.I(\beepboop.inst.counter[6] ),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1765_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1766_ (.A1(_1295_),
    .A2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1767_ (.A1(_1294_),
    .A2(_1298_),
    .B(_1270_),
    .C(_1272_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1768_ (.A1(_1280_),
    .A2(_1299_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1769_ (.A1(_1289_),
    .A2(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1770_ (.I(_1300_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1771_ (.A1(_1276_),
    .A2(_1273_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1772_ (.A1(_1292_),
    .A2(_1301_),
    .B(_1290_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1773_ (.I(\beepboop.inst.counter[10] ),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1774_ (.I(\beepboop.inst.counter[8] ),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1775_ (.A1(_1303_),
    .A2(_1304_),
    .A3(_1295_),
    .A4(_1296_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1776_ (.I(\beepboop.inst.counter[9] ),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1777_ (.A1(_1303_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1778_ (.A1(_1302_),
    .A2(_1305_),
    .B(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1779_ (.A1(\beepboop.inst.counter[10] ),
    .A2(\beepboop.inst.counter[9] ),
    .A3(_1277_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1780_ (.A1(\beepboop.inst.counter[3] ),
    .A2(_1273_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1781_ (.A1(_1279_),
    .A2(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1782_ (.A1(_1292_),
    .A2(_1311_),
    .B(_1290_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1783_ (.A1(_1309_),
    .A2(_1312_),
    .B(_1270_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(_1272_),
    .A2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1785_ (.A1(_1308_),
    .A2(_1314_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1786_ (.A1(\beepboop.inst.counter[10] ),
    .A2(_1306_),
    .A3(\beepboop.inst.counter[8] ),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1787_ (.I(_1284_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1788_ (.A1(\beepboop.inst.counter[3] ),
    .A2(\beepboop.inst.counter[2] ),
    .B(_1275_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1789_ (.I(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1790_ (.A1(_1290_),
    .A2(\beepboop.inst.counter[4] ),
    .B(_1318_),
    .C(_1296_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1791_ (.A1(_1316_),
    .A2(_1319_),
    .B(_1277_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1792_ (.A1(_1278_),
    .A2(_1315_),
    .B1(_1320_),
    .B2(_1304_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1793_ (.A1(_1306_),
    .A2(_1321_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1794_ (.A1(_1291_),
    .A2(_1293_),
    .B(_1295_),
    .C(_1297_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1795_ (.A1(_1292_),
    .A2(_1301_),
    .B(_1296_),
    .C(_1291_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1796_ (.A1(_1316_),
    .A2(_1324_),
    .B(_1315_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1797_ (.A1(_1308_),
    .A2(_1322_),
    .B1(_1323_),
    .B2(_1325_),
    .C(_1314_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1798_ (.A1(_1293_),
    .A2(_1318_),
    .B(_1277_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1799_ (.A1(\beepboop.inst.counter[11] ),
    .A2(_1270_),
    .A3(_1282_),
    .A4(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1800_ (.A1(_1326_),
    .A2(_1328_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1801_ (.I(\ttA_0.io_out[0] ),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1802_ (.I(_1329_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1803_ (.I(_1330_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1804_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1805_ (.I(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1806_ (.I(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1807_ (.I(net9),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1808_ (.I(net10),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1809_ (.A1(_1335_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1810_ (.I(net11),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1811_ (.A1(_1338_),
    .A2(net10),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1812_ (.A1(_1338_),
    .A2(net9),
    .A3(_1336_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1813_ (.A1(_1337_),
    .A2(_1339_),
    .A3(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1814_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1815_ (.I(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1816_ (.A1(\ttA_6.counter[15] ),
    .A2(\ttA_6.counter[14] ),
    .A3(\ttA_6.counter[13] ),
    .A4(\ttA_6.counter[12] ),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1817_ (.I(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1818_ (.I(\ttA_6.counter[11] ),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1819_ (.I(\ttA_6.counter[7] ),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1820_ (.I(\ttA_6.counter[4] ),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1821_ (.I(\ttA_6.counter[6] ),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1822_ (.I(\ttA_6.counter[5] ),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1823_ (.I(_1350_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1824_ (.A1(_1348_),
    .A2(\ttA_6.counter[3] ),
    .B(_1349_),
    .C(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1825_ (.A1(\ttA_6.counter[10] ),
    .A2(\ttA_6.counter[9] ),
    .A3(\ttA_6.counter[8] ),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1826_ (.A1(_1347_),
    .A2(_1352_),
    .B(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1827_ (.A1(_1346_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1828_ (.A1(_1345_),
    .A2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1829_ (.A1(\ttA_6.counter[7] ),
    .A2(_1349_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1830_ (.I(\ttA_6.counter[3] ),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1831_ (.A1(_1351_),
    .A2(_1348_),
    .A3(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1832_ (.I(_1353_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1833_ (.A1(\ttA_6.counter[11] ),
    .A2(_1344_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1834_ (.A1(_1357_),
    .A2(_1359_),
    .B(_1360_),
    .C(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1835_ (.A1(_1338_),
    .A2(_1335_),
    .A3(_1336_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1836_ (.I(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(_1362_),
    .A2(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1838_ (.A1(net9),
    .A2(_1339_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1839_ (.I(_1366_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1840_ (.I(_1076_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1841_ (.I(net32),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1842_ (.I(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1843_ (.A1(_1370_),
    .A2(net95),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1844_ (.I(net32),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1845_ (.I(net95),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1846_ (.A1(_1372_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1847_ (.A1(_1374_),
    .A2(_1371_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1848_ (.A1(_1142_),
    .A2(_1076_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1849_ (.I(_1372_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1850_ (.A1(_1377_),
    .A2(_1373_),
    .B(_1166_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1851_ (.A1(_1368_),
    .A2(_1371_),
    .B1(_1375_),
    .B2(_1376_),
    .C(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1852_ (.A1(_1338_),
    .A2(_1335_),
    .A3(net10),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1853_ (.A1(net11),
    .A2(_1335_),
    .A3(_1336_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1854_ (.A1(\ttA_4.pwm_signal ),
    .A2(_1380_),
    .B1(_1381_),
    .B2(\ttA_2.io_out[0] ),
    .C(_1341_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1855_ (.A1(_1356_),
    .A2(_1365_),
    .B1(_1367_),
    .B2(_1379_),
    .C(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1856_ (.I(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1857_ (.A1(_1334_),
    .A2(_1343_),
    .B(_1384_),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1858_ (.I(\ttA_6.counter[2] ),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1859_ (.I(\ttA_6.counter[0] ),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1860_ (.I(\ttA_6.counter[7] ),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1861_ (.A1(_1387_),
    .A2(_1349_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1862_ (.A1(_1359_),
    .A2(_1388_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1863_ (.A1(_1385_),
    .A2(\ttA_6.counter[1] ),
    .A3(_1386_),
    .A4(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1864_ (.I(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1865_ (.A1(_1364_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1866_ (.I(\ttA_0.io_out[1] ),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1867_ (.I(_1393_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1868_ (.I(_1394_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1869_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1870_ (.I(_1342_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1871_ (.I(_1381_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1872_ (.I(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1873_ (.I(_1366_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1874_ (.I(_1370_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1875_ (.A1(_1127_),
    .A2(_1076_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1876_ (.I(net95),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1877_ (.A1(_1168_),
    .A2(_1078_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1878_ (.A1(_1403_),
    .A2(_1376_),
    .A3(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1879_ (.A1(_1077_),
    .A2(net32),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1880_ (.A1(net3),
    .A2(_1369_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1881_ (.I(_1406_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1882_ (.A1(_1373_),
    .A2(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1883_ (.A1(_1168_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1884_ (.A1(_1403_),
    .A2(_1406_),
    .B1(_1407_),
    .B2(_1410_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1885_ (.A1(_1401_),
    .A2(_1402_),
    .B(_1405_),
    .C(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1886_ (.A1(_1400_),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1887_ (.A1(_1396_),
    .A2(_1397_),
    .B1(_1399_),
    .B2(_1130_),
    .C(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1888_ (.A1(_1362_),
    .A2(_1392_),
    .B(_1414_),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1889_ (.A1(_1376_),
    .A2(_1375_),
    .A3(_1405_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1890_ (.I(\ttA_0.io_out[2] ),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1891_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1892_ (.I(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1893_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1894_ (.I(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1895_ (.A1(_1420_),
    .A2(_1397_),
    .B1(_1399_),
    .B2(_1134_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1896_ (.A1(_1360_),
    .A2(_1361_),
    .A3(_1390_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1897_ (.A1(_1356_),
    .A2(_1422_),
    .B(_1364_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1898_ (.A1(_1367_),
    .A2(_1415_),
    .B(_1421_),
    .C(_1423_),
    .ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1899_ (.I(_1078_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1900_ (.A1(_1406_),
    .A2(_1407_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1901_ (.I(_1129_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1902_ (.A1(_0003_),
    .A2(_1403_),
    .B1(_1424_),
    .B2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1903_ (.A1(_1149_),
    .A2(_1371_),
    .A3(_1409_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1904_ (.A1(_1426_),
    .A2(_1427_),
    .B(_1367_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1905_ (.A1(\ttA_2.io_out[3] ),
    .A2(_1399_),
    .B(_1428_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1906_ (.I(_1340_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1907_ (.I(\ttA_0.io_out[3] ),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1908_ (.I(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1909_ (.I(_1432_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1910_ (.I(_1433_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1911_ (.I(\ttA_6.counter[10] ),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1912_ (.I(\ttA_6.counter[8] ),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1913_ (.A1(\ttA_6.counter[3] ),
    .A2(\ttA_6.counter[2] ),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1914_ (.I(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1915_ (.A1(_1348_),
    .A2(_1438_),
    .B(_1350_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1916_ (.A1(_1357_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1917_ (.I(\ttA_6.counter[9] ),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1918_ (.A1(_1436_),
    .A2(_1440_),
    .B(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1919_ (.A1(_1435_),
    .A2(_1442_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1920_ (.A1(_1346_),
    .A2(_1360_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1921_ (.A1(_1363_),
    .A2(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1922_ (.A1(\ttA_6.counter[1] ),
    .A2(_1386_),
    .B(_1438_),
    .C(_1351_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1923_ (.I(_1350_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1924_ (.I(\ttA_6.counter[4] ),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1925_ (.A1(_1447_),
    .A2(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1926_ (.I(\ttA_6.counter[8] ),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1927_ (.A1(\ttA_6.counter[11] ),
    .A2(\ttA_6.counter[10] ),
    .A3(\ttA_6.counter[9] ),
    .A4(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1928_ (.A1(_1388_),
    .A2(_1446_),
    .A3(_1449_),
    .A4(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(_1345_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1930_ (.A1(_1443_),
    .A2(_1445_),
    .A3(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1931_ (.A1(_1220_),
    .A2(_1430_),
    .B1(_1343_),
    .B2(_1434_),
    .C(_1454_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1932_ (.A1(_1429_),
    .A2(_1455_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(\ttA_6.counter[6] ),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1934_ (.A1(_1456_),
    .A2(_1448_),
    .A3(_1358_),
    .A4(\ttA_6.counter[2] ),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1935_ (.A1(_1456_),
    .A2(_1447_),
    .B(_1387_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1936_ (.A1(_1387_),
    .A2(_1456_),
    .B1(_1457_),
    .B2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1937_ (.A1(_1351_),
    .A2(_1348_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1938_ (.A1(\ttA_6.counter[4] ),
    .A2(_1438_),
    .B(_1349_),
    .C(_1350_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1939_ (.A1(_1347_),
    .A2(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1940_ (.A1(_1357_),
    .A2(_1460_),
    .B(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1941_ (.A1(_1441_),
    .A2(_1436_),
    .A3(_1389_),
    .A4(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1942_ (.A1(_1436_),
    .A2(_1459_),
    .B(_1464_),
    .C(_1443_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1943_ (.A1(_1358_),
    .A2(_1385_),
    .B(_1447_),
    .C(_1448_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1944_ (.A1(_1346_),
    .A2(_1360_),
    .A3(_1388_),
    .A4(_1466_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1945_ (.A1(_1444_),
    .A2(_1465_),
    .B(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1946_ (.A1(_1453_),
    .A2(_1468_),
    .B(_1364_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1947_ (.I(\ttA_0.io_out[4] ),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1948_ (.I(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1949_ (.A1(_1078_),
    .A2(_1401_),
    .B(_1373_),
    .C(_1400_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1950_ (.A1(\ttA_2.io_out[4] ),
    .A2(_1398_),
    .B(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1951_ (.A1(_1425_),
    .A2(_1400_),
    .A3(_1408_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1952_ (.A1(_1243_),
    .A2(_1430_),
    .B1(_1397_),
    .B2(_1471_),
    .C(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1953_ (.A1(_1469_),
    .A2(_1475_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1954_ (.I(\ttA_0.io_out[5] ),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1955_ (.I(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1956_ (.I(_1234_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1957_ (.I(\ttA_1.top.backend.rptr[1] ),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1958_ (.I0(\ttA_1.top.data[4][0] ),
    .I1(\ttA_1.top.data[5][0] ),
    .I2(\ttA_1.top.data[6][0] ),
    .I3(\ttA_1.top.data[7][0] ),
    .S0(_1478_),
    .S1(_1479_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1959_ (.I(_1234_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1960_ (.I(\ttA_1.top.data[1][0] ),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1961_ (.A1(_1481_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1962_ (.A1(_1252_),
    .A2(\ttA_1.top.data[0][0] ),
    .B(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1963_ (.I(\ttA_1.top.data[3][0] ),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1964_ (.A1(_1478_),
    .A2(_1485_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1965_ (.A1(_1235_),
    .A2(\ttA_1.top.data[2][0] ),
    .B(_1486_),
    .C(_1233_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1966_ (.A1(_1250_),
    .A2(_1484_),
    .B(_1487_),
    .C(_1231_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1967_ (.A1(_1248_),
    .A2(_1480_),
    .B(_1488_),
    .C(_1430_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1968_ (.A1(_1144_),
    .A2(_1398_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1969_ (.A1(_1367_),
    .A2(_1411_),
    .B(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1970_ (.A1(_1397_),
    .A2(_1454_),
    .A3(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1971_ (.A1(_1477_),
    .A2(_1343_),
    .B1(_1489_),
    .B2(_1492_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1972_ (.I0(\ttA_1.top.data[2][1] ),
    .I1(\ttA_1.top.data[3][1] ),
    .S(_1481_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1973_ (.I(\ttA_1.top.data[1][1] ),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1974_ (.A1(_1235_),
    .A2(\ttA_1.top.data[0][1] ),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1975_ (.A1(_1252_),
    .A2(_1494_),
    .B(_1495_),
    .C(_1479_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1976_ (.A1(_1250_),
    .A2(_1493_),
    .B(_1496_),
    .C(\ttA_1.top.backend.rptr[2] ),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1977_ (.I0(\ttA_1.top.data[4][1] ),
    .I1(\ttA_1.top.data[5][1] ),
    .I2(\ttA_1.top.data[6][1] ),
    .I3(\ttA_1.top.data[7][1] ),
    .S0(_1481_),
    .S1(_1479_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1978_ (.A1(_1248_),
    .A2(_1498_),
    .B(_1430_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1979_ (.I(\ttA_0.io_out[6] ),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1980_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1981_ (.I(_1501_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1982_ (.A1(_1149_),
    .A2(_1377_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1983_ (.I(_1407_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1984_ (.A1(_1403_),
    .A2(_1503_),
    .B(_1404_),
    .C(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1985_ (.A1(_1409_),
    .A2(_1505_),
    .B(_1400_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1986_ (.A1(_1502_),
    .A2(_1342_),
    .B1(_1398_),
    .B2(_1147_),
    .C(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1987_ (.A1(_1497_),
    .A2(_1499_),
    .B(_1507_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1988_ (.I(\ttA_0.io_out[7] ),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1989_ (.I(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1990_ (.I0(\ttA_1.top.data[4][2] ),
    .I1(\ttA_1.top.data[5][2] ),
    .I2(\ttA_1.top.data[6][2] ),
    .I3(\ttA_1.top.data[7][2] ),
    .S0(_1478_),
    .S1(_1479_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1991_ (.I(\ttA_1.top.data[1][2] ),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1992_ (.A1(_1481_),
    .A2(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1993_ (.A1(_1252_),
    .A2(\ttA_1.top.data[0][2] ),
    .B(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1994_ (.I(\ttA_1.top.data[3][2] ),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1995_ (.A1(_1478_),
    .A2(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1996_ (.A1(_1235_),
    .A2(\ttA_1.top.data[2][2] ),
    .B(_1515_),
    .C(_1233_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1997_ (.A1(_1250_),
    .A2(_1513_),
    .B(_1516_),
    .C(_1231_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1998_ (.A1(_1248_),
    .A2(_1510_),
    .B(_1517_),
    .C(_1340_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1999_ (.A1(\ttA_2.io_out[7] ),
    .A2(_1399_),
    .B(_1472_),
    .C(_1342_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2000_ (.A1(_1509_),
    .A2(_1343_),
    .B1(_1518_),
    .B2(_1519_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2001_ (.I(\ttA_0.io_out[3] ),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2002_ (.I(_1520_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2003_ (.I(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2004_ (.I(\ttA_0.io_out[2] ),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2005_ (.I(\ttA_0.io_out[0] ),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2006_ (.I(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2007_ (.I0(\ttA_0.prog[8][2] ),
    .I1(\ttA_0.prog[9][2] ),
    .I2(\ttA_0.prog[10][2] ),
    .I3(\ttA_0.prog[11][2] ),
    .S0(_0259_),
    .S1(_1393_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2008_ (.A1(_0257_),
    .A2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2009_ (.I(\ttA_0.io_out[2] ),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2010_ (.I(_0262_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2011_ (.I0(\ttA_0.prog[12][2] ),
    .I1(\ttA_0.prog[13][2] ),
    .I2(\ttA_0.prog[14][2] ),
    .I3(\ttA_0.prog[15][2] ),
    .S0(_0259_),
    .S1(_1393_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2012_ (.A1(_0263_),
    .A2(_0264_),
    .B(_1431_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2013_ (.I(\ttA_0.io_out[0] ),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2014_ (.I(\ttA_0.io_out[1] ),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2015_ (.I(_0267_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2016_ (.I0(\ttA_0.prog[0][2] ),
    .I1(\ttA_0.prog[1][2] ),
    .I2(\ttA_0.prog[2][2] ),
    .I3(\ttA_0.prog[3][2] ),
    .S0(_0266_),
    .S1(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2017_ (.A1(_1416_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2018_ (.I0(\ttA_0.prog[4][2] ),
    .I1(\ttA_0.prog[5][2] ),
    .I2(\ttA_0.prog[6][2] ),
    .I3(\ttA_0.prog[7][2] ),
    .S0(_0259_),
    .S1(_1393_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2019_ (.A1(_0263_),
    .A2(_0271_),
    .B(_1520_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2020_ (.A1(_0261_),
    .A2(_0265_),
    .B1(_0270_),
    .B2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2021_ (.I(\ttA_0.io_out[1] ),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2022_ (.I0(\ttA_0.prog[0][3] ),
    .I1(\ttA_0.prog[1][3] ),
    .I2(\ttA_0.prog[2][3] ),
    .I3(\ttA_0.prog[3][3] ),
    .S0(_0258_),
    .S1(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2023_ (.A1(_1416_),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2024_ (.I0(\ttA_0.prog[4][3] ),
    .I1(\ttA_0.prog[5][3] ),
    .I2(\ttA_0.prog[6][3] ),
    .I3(\ttA_0.prog[7][3] ),
    .S0(_0266_),
    .S1(_0274_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2025_ (.A1(_0262_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2026_ (.I0(\ttA_0.prog[8][3] ),
    .I1(\ttA_0.prog[9][3] ),
    .I2(\ttA_0.prog[10][3] ),
    .I3(\ttA_0.prog[11][3] ),
    .S0(_0266_),
    .S1(_0268_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2027_ (.A1(_1416_),
    .A2(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2028_ (.I0(\ttA_0.prog[12][3] ),
    .I1(\ttA_0.prog[13][3] ),
    .I2(\ttA_0.prog[14][3] ),
    .I3(\ttA_0.prog[15][3] ),
    .S0(_0266_),
    .S1(_0268_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2029_ (.A1(_0263_),
    .A2(_0281_),
    .B(_1431_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2030_ (.A1(_1433_),
    .A2(_0276_),
    .A3(_0278_),
    .B1(_0280_),
    .B2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2031_ (.A1(_0273_),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2032_ (.I0(\ttA_0.prog[8][0] ),
    .I1(\ttA_0.prog[9][0] ),
    .I2(\ttA_0.prog[10][0] ),
    .I3(\ttA_0.prog[11][0] ),
    .S0(_1330_),
    .S1(_1394_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2033_ (.A1(_1417_),
    .A2(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2034_ (.I(_0263_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2035_ (.I0(\ttA_0.prog[12][0] ),
    .I1(\ttA_0.prog[13][0] ),
    .I2(\ttA_0.prog[14][0] ),
    .I3(\ttA_0.prog[15][0] ),
    .S0(_1330_),
    .S1(_1394_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2036_ (.I(_1431_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2037_ (.A1(_0287_),
    .A2(_0288_),
    .B(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2038_ (.A1(_0286_),
    .A2(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2039_ (.I(\ttA_0.io_out[2] ),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2040_ (.I(_0259_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2041_ (.I(_0267_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2042_ (.I0(\ttA_0.prog[0][0] ),
    .I1(\ttA_0.prog[1][0] ),
    .I2(\ttA_0.prog[2][0] ),
    .I3(\ttA_0.prog[3][0] ),
    .S0(_0293_),
    .S1(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2043_ (.A1(_0292_),
    .A2(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2044_ (.I(_0262_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2045_ (.I(_1329_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2046_ (.I(_0274_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2047_ (.I0(\ttA_0.prog[4][0] ),
    .I1(\ttA_0.prog[5][0] ),
    .I2(\ttA_0.prog[6][0] ),
    .I3(\ttA_0.prog[7][0] ),
    .S0(_0298_),
    .S1(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2048_ (.A1(_0297_),
    .A2(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2049_ (.A1(_1433_),
    .A2(_0296_),
    .A3(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2050_ (.I0(\ttA_0.prog[8][1] ),
    .I1(\ttA_0.prog[9][1] ),
    .I2(\ttA_0.prog[10][1] ),
    .I3(\ttA_0.prog[11][1] ),
    .S0(_0298_),
    .S1(_0299_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2051_ (.A1(_1417_),
    .A2(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2052_ (.I0(\ttA_0.prog[12][1] ),
    .I1(\ttA_0.prog[13][1] ),
    .I2(\ttA_0.prog[14][1] ),
    .I3(\ttA_0.prog[15][1] ),
    .S0(_0298_),
    .S1(_0299_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2053_ (.A1(_0287_),
    .A2(_0305_),
    .B(_0289_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2054_ (.I0(\ttA_0.prog[0][1] ),
    .I1(\ttA_0.prog[1][1] ),
    .I2(\ttA_0.prog[2][1] ),
    .I3(\ttA_0.prog[3][1] ),
    .S0(_0293_),
    .S1(_0294_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2055_ (.A1(_1417_),
    .A2(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2056_ (.I0(\ttA_0.prog[4][1] ),
    .I1(\ttA_0.prog[5][1] ),
    .I2(\ttA_0.prog[6][1] ),
    .I3(\ttA_0.prog[7][1] ),
    .S0(_0298_),
    .S1(_0299_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2057_ (.A1(_0297_),
    .A2(_0309_),
    .B(_0255_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2058_ (.A1(_0304_),
    .A2(_0306_),
    .B1(_0308_),
    .B2(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2059_ (.A1(_0291_),
    .A2(_0302_),
    .B(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2060_ (.A1(_1091_),
    .A2(_1504_),
    .A3(_0284_),
    .A4(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2061_ (.I(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2062_ (.I(_0313_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2063_ (.I0(\ttA_0.data[8][3] ),
    .I1(\ttA_0.data[9][3] ),
    .I2(\ttA_0.data[10][3] ),
    .I3(\ttA_0.data[11][3] ),
    .S0(_1331_),
    .S1(_1395_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2064_ (.A1(_1418_),
    .A2(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2065_ (.I(_0287_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2066_ (.I0(\ttA_0.data[12][3] ),
    .I1(\ttA_0.data[14][3] ),
    .I2(\ttA_0.data[13][3] ),
    .I3(\ttA_0.data[15][3] ),
    .S0(_1395_),
    .S1(_1331_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2067_ (.A1(_0318_),
    .A2(_0319_),
    .B(_1434_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2068_ (.I0(\ttA_0.data[4][3] ),
    .I1(\ttA_0.data[6][3] ),
    .I2(\ttA_0.data[5][3] ),
    .I3(\ttA_0.data[7][3] ),
    .S0(_1395_),
    .S1(_1331_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2069_ (.I0(\ttA_0.data[0][3] ),
    .I1(\ttA_0.data[1][3] ),
    .I2(\ttA_0.data[2][3] ),
    .I3(\ttA_0.data[3][3] ),
    .S0(_1330_),
    .S1(_1394_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2070_ (.A1(_1418_),
    .A2(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2071_ (.A1(_0287_),
    .A2(_0321_),
    .B(_0323_),
    .C(_0256_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2072_ (.A1(_0317_),
    .A2(_0320_),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2073_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2074_ (.A1(_0315_),
    .A2(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2075_ (.A1(_0256_),
    .A2(_0314_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2076_ (.I(_0258_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2077_ (.I(_0267_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2078_ (.I0(\ttA_0.data[0][2] ),
    .I1(\ttA_0.data[1][2] ),
    .I2(\ttA_0.data[2][2] ),
    .I3(\ttA_0.data[3][2] ),
    .S0(_0329_),
    .S1(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2079_ (.A1(_0257_),
    .A2(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2080_ (.I(_0262_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2081_ (.I(_0267_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2082_ (.I(_0258_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2083_ (.I0(\ttA_0.data[4][2] ),
    .I1(\ttA_0.data[6][2] ),
    .I2(\ttA_0.data[5][2] ),
    .I3(\ttA_0.data[7][2] ),
    .S0(_0334_),
    .S1(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2084_ (.A1(_0333_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2085_ (.I0(\ttA_0.data[8][2] ),
    .I1(\ttA_0.data[9][2] ),
    .I2(\ttA_0.data[10][2] ),
    .I3(\ttA_0.data[11][2] ),
    .S0(_0329_),
    .S1(_0294_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2086_ (.A1(_0292_),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2087_ (.I0(\ttA_0.data[12][2] ),
    .I1(\ttA_0.data[14][2] ),
    .I2(\ttA_0.data[13][2] ),
    .I3(\ttA_0.data[15][2] ),
    .S0(_0334_),
    .S1(_0335_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2088_ (.A1(_0333_),
    .A2(_0340_),
    .B(_0289_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2089_ (.A1(_0289_),
    .A2(_0332_),
    .A3(_0337_),
    .B1(_0339_),
    .B2(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2090_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2091_ (.I(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2092_ (.I(_0313_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2093_ (.A1(_1418_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2094_ (.A1(_0314_),
    .A2(_0344_),
    .B(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2095_ (.A1(_0328_),
    .A2(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2096_ (.A1(_1127_),
    .A2(_1407_),
    .B(_0314_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2097_ (.I(_0315_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2098_ (.I0(\ttA_0.data[0][0] ),
    .I1(\ttA_0.data[1][0] ),
    .I2(\ttA_0.data[2][0] ),
    .I3(\ttA_0.data[3][0] ),
    .S0(_0329_),
    .S1(_0294_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2099_ (.A1(_0292_),
    .A2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2100_ (.I0(\ttA_0.data[4][0] ),
    .I1(\ttA_0.data[6][0] ),
    .I2(\ttA_0.data[5][0] ),
    .I3(\ttA_0.data[7][0] ),
    .S0(_0330_),
    .S1(_0293_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2101_ (.A1(_0297_),
    .A2(_0353_),
    .B(_0255_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2102_ (.I0(\ttA_0.data[8][0] ),
    .I1(\ttA_0.data[9][0] ),
    .I2(\ttA_0.data[10][0] ),
    .I3(\ttA_0.data[11][0] ),
    .S0(_0329_),
    .S1(_0330_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2103_ (.A1(_0292_),
    .A2(_0355_),
    .B(_1432_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2104_ (.I0(\ttA_0.data[12][0] ),
    .I1(\ttA_0.data[14][0] ),
    .I2(\ttA_0.data[13][0] ),
    .I3(\ttA_0.data[15][0] ),
    .S0(_0330_),
    .S1(_0293_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2105_ (.A1(_0297_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2106_ (.A1(_0352_),
    .A2(_0354_),
    .B1(_0356_),
    .B2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2107_ (.I(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2108_ (.I(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2109_ (.I(_0361_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2110_ (.A1(_1332_),
    .A2(_0345_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2111_ (.A1(_0350_),
    .A2(_0362_),
    .B(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2112_ (.I0(\ttA_0.data[8][1] ),
    .I1(\ttA_0.data[9][1] ),
    .I2(\ttA_0.data[10][1] ),
    .I3(\ttA_0.data[11][1] ),
    .S0(_1329_),
    .S1(_0334_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2113_ (.A1(_0257_),
    .A2(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2114_ (.I0(\ttA_0.data[12][1] ),
    .I1(\ttA_0.data[14][1] ),
    .I2(\ttA_0.data[13][1] ),
    .I3(\ttA_0.data[15][1] ),
    .S0(_0268_),
    .S1(_0335_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2115_ (.A1(_0333_),
    .A2(_0367_),
    .B(_1432_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2116_ (.I0(\ttA_0.data[0][1] ),
    .I1(\ttA_0.data[1][1] ),
    .I2(\ttA_0.data[2][1] ),
    .I3(\ttA_0.data[3][1] ),
    .S0(_1329_),
    .S1(_0334_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2117_ (.A1(_0257_),
    .A2(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2118_ (.I0(\ttA_0.data[4][1] ),
    .I1(\ttA_0.data[6][1] ),
    .I2(\ttA_0.data[5][1] ),
    .I3(\ttA_0.data[7][1] ),
    .S0(_0274_),
    .S1(_0335_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2119_ (.A1(_0333_),
    .A2(_0371_),
    .B(_0255_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2120_ (.A1(_0366_),
    .A2(_0368_),
    .B1(_0370_),
    .B2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2121_ (.I(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2122_ (.A1(_0315_),
    .A2(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2123_ (.I(_1396_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2124_ (.A1(_0376_),
    .A2(_0315_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2125_ (.A1(_0375_),
    .A2(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2126_ (.A1(_0349_),
    .A2(_0364_),
    .A3(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2127_ (.A1(_0348_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2128_ (.I(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2129_ (.I(_0350_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2130_ (.I(_0350_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(_1126_),
    .A2(_0383_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2132_ (.A1(_1471_),
    .A2(_0382_),
    .B(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2133_ (.I(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2134_ (.I(_0380_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2135_ (.A1(\ttA_0.data[1][0] ),
    .A2(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2136_ (.I(_1372_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2137_ (.I(_0389_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2138_ (.A1(_0381_),
    .A2(_0386_),
    .B(_0388_),
    .C(_0390_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2139_ (.I(_1476_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2140_ (.I(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2141_ (.A1(_1153_),
    .A2(_0383_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2142_ (.A1(_0392_),
    .A2(_0382_),
    .B(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2143_ (.I(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2144_ (.A1(\ttA_0.data[1][1] ),
    .A2(_0387_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2145_ (.A1(_0381_),
    .A2(_0395_),
    .B(_0396_),
    .C(_0390_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2146_ (.I(_1083_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2147_ (.A1(_0397_),
    .A2(_0383_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2148_ (.A1(_1502_),
    .A2(_0382_),
    .B(_0398_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2149_ (.I(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2150_ (.A1(\ttA_0.data[1][2] ),
    .A2(_0387_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2151_ (.A1(_0381_),
    .A2(_0400_),
    .B(_0401_),
    .C(_0390_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2152_ (.I(_1508_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2153_ (.A1(_1159_),
    .A2(_0383_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2154_ (.A1(_0402_),
    .A2(_0382_),
    .B(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2155_ (.I(_0404_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2156_ (.A1(\ttA_0.data[1][3] ),
    .A2(_0387_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2157_ (.I(_1377_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2158_ (.I(_0407_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2159_ (.A1(_0381_),
    .A2(_0405_),
    .B(_0406_),
    .C(_0408_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2160_ (.I(_0359_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2161_ (.A1(_1333_),
    .A2(_0345_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2162_ (.A1(_0350_),
    .A2(_0409_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2163_ (.A1(_0349_),
    .A2(_0411_),
    .A3(_0378_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2164_ (.A1(_0348_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2165_ (.I(_0413_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2166_ (.I(_0413_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2167_ (.A1(\ttA_0.data[0][0] ),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2168_ (.A1(_0386_),
    .A2(_0414_),
    .B(_0416_),
    .C(_0408_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2169_ (.A1(\ttA_0.data[0][1] ),
    .A2(_0415_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2170_ (.A1(_0395_),
    .A2(_0414_),
    .B(_0417_),
    .C(_0408_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2171_ (.A1(\ttA_0.data[0][2] ),
    .A2(_0415_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2172_ (.A1(_0400_),
    .A2(_0414_),
    .B(_0418_),
    .C(_0408_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2173_ (.A1(\ttA_0.data[0][3] ),
    .A2(_0415_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2174_ (.I(_1372_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2175_ (.I(_0420_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2176_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2177_ (.A1(_0405_),
    .A2(_0414_),
    .B(_0419_),
    .C(_0422_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2178_ (.I(_1197_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2179_ (.A1(_1143_),
    .A2(\ttA_1.top.frontend.wptr[0] ),
    .A3(_1220_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2180_ (.A1(_1225_),
    .A2(_1209_),
    .A3(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2181_ (.I(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2182_ (.A1(\ttA_1.top.data[6][0] ),
    .A2(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2183_ (.A1(_0423_),
    .A2(_0426_),
    .B(_0427_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2184_ (.I(_0397_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(\ttA_1.top.data[6][1] ),
    .A2(_0425_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2186_ (.A1(_0428_),
    .A2(_0426_),
    .B(_0429_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2187_ (.I(_1180_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(\ttA_1.top.data[6][2] ),
    .A2(_0425_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2189_ (.A1(_0430_),
    .A2(_0426_),
    .B(_0431_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2190_ (.I(_1197_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2191_ (.I(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2192_ (.A1(_1208_),
    .A2(_1228_),
    .A3(_1222_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2193_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2194_ (.A1(\ttA_1.top.data[5][0] ),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2195_ (.A1(_0433_),
    .A2(_0435_),
    .B(_0436_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2196_ (.I(_0397_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2197_ (.I(_0437_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2198_ (.A1(\ttA_1.top.data[5][1] ),
    .A2(_0434_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2199_ (.A1(_0438_),
    .A2(_0435_),
    .B(_0439_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2200_ (.I(_1160_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2201_ (.A1(\ttA_1.top.data[5][2] ),
    .A2(_0434_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2202_ (.A1(_0440_),
    .A2(_0435_),
    .B(_0441_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2203_ (.I(_1197_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2204_ (.A1(_1225_),
    .A2(_1228_),
    .A3(_0424_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2205_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2206_ (.A1(\ttA_1.top.data[4][0] ),
    .A2(_0444_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2207_ (.A1(_0442_),
    .A2(_0444_),
    .B(_0445_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2208_ (.I(_0397_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2209_ (.A1(\ttA_1.top.data[4][1] ),
    .A2(_0443_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2210_ (.A1(_0446_),
    .A2(_0444_),
    .B(_0447_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2211_ (.I(_1160_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2212_ (.A1(\ttA_1.top.data[4][2] ),
    .A2(_0443_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2213_ (.A1(_0448_),
    .A2(_0444_),
    .B(_0449_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2214_ (.A1(_1225_),
    .A2(_1226_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2215_ (.I(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_1123_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2217_ (.A1(_0452_),
    .A2(_0451_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2218_ (.A1(_1485_),
    .A2(_0451_),
    .B(_0453_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2219_ (.A1(\ttA_1.top.data[3][1] ),
    .A2(_0450_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2220_ (.A1(_0438_),
    .A2(_0451_),
    .B(_0454_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2221_ (.A1(_1196_),
    .A2(_0450_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2222_ (.A1(_1514_),
    .A2(_0451_),
    .B(_0455_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2223_ (.A1(_1208_),
    .A2(_1228_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2224_ (.A1(_0456_),
    .A2(_0424_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2225_ (.I(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2226_ (.A1(\ttA_1.top.data[2][0] ),
    .A2(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2227_ (.A1(_0442_),
    .A2(_0458_),
    .B(_0459_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2228_ (.A1(\ttA_1.top.data[2][1] ),
    .A2(_0457_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2229_ (.A1(_0446_),
    .A2(_0458_),
    .B(_0460_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2230_ (.A1(\ttA_1.top.data[2][2] ),
    .A2(_0457_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2231_ (.A1(_0448_),
    .A2(_0458_),
    .B(_0461_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2232_ (.A1(_1208_),
    .A2(_1209_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(_1222_),
    .A2(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2234_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2235_ (.A1(\ttA_1.top.data[1][0] ),
    .A2(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2236_ (.A1(_0442_),
    .A2(_0464_),
    .B(_0465_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2237_ (.A1(\ttA_1.top.data[1][1] ),
    .A2(_0463_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2238_ (.A1(_0446_),
    .A2(_0464_),
    .B(_0466_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2239_ (.A1(\ttA_1.top.data[1][2] ),
    .A2(_0463_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2240_ (.A1(_0448_),
    .A2(_0464_),
    .B(_0467_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2241_ (.A1(_0424_),
    .A2(_0462_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2242_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2243_ (.A1(\ttA_1.top.data[0][0] ),
    .A2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2244_ (.A1(_0442_),
    .A2(_0469_),
    .B(_0470_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2245_ (.A1(\ttA_1.top.data[0][1] ),
    .A2(_0468_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2246_ (.A1(_0446_),
    .A2(_0469_),
    .B(_0471_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2247_ (.A1(\ttA_1.top.data[0][2] ),
    .A2(_0468_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2248_ (.A1(_0448_),
    .A2(_0469_),
    .B(_0472_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2249_ (.I(_0343_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_0318_),
    .A2(_0345_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2251_ (.A1(_0314_),
    .A2(_0473_),
    .B(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2252_ (.A1(_0328_),
    .A2(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2253_ (.A1(_0379_),
    .A2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2254_ (.I(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2255_ (.I(_0477_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2256_ (.A1(\ttA_0.data[9][0] ),
    .A2(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2257_ (.A1(_0386_),
    .A2(_0478_),
    .B(_0480_),
    .C(_0422_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2258_ (.A1(\ttA_0.data[9][1] ),
    .A2(_0479_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2259_ (.A1(_0395_),
    .A2(_0478_),
    .B(_0481_),
    .C(_0422_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2260_ (.A1(\ttA_0.data[9][2] ),
    .A2(_0479_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2261_ (.A1(_0400_),
    .A2(_0478_),
    .B(_0482_),
    .C(_0422_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(\ttA_0.data[9][3] ),
    .A2(_0479_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2263_ (.I(_0421_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2264_ (.A1(_0405_),
    .A2(_0478_),
    .B(_0483_),
    .C(_0484_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2265_ (.A1(_0349_),
    .A2(_0364_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2266_ (.I(_0378_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2267_ (.A1(_0328_),
    .A2(_0475_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2268_ (.A1(_0485_),
    .A2(_0486_),
    .A3(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2269_ (.I(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2270_ (.I(_0488_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2271_ (.A1(\ttA_0.data[7][0] ),
    .A2(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2272_ (.A1(_0386_),
    .A2(_0489_),
    .B(_0491_),
    .C(_0484_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2273_ (.A1(\ttA_0.data[7][1] ),
    .A2(_0490_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2274_ (.A1(_0395_),
    .A2(_0489_),
    .B(_0492_),
    .C(_0484_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2275_ (.A1(\ttA_0.data[7][2] ),
    .A2(_0490_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2276_ (.A1(_0400_),
    .A2(_0489_),
    .B(_0493_),
    .C(_0484_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2277_ (.A1(\ttA_0.data[7][3] ),
    .A2(_0490_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2278_ (.I(_0421_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2279_ (.A1(_0405_),
    .A2(_0489_),
    .B(_0494_),
    .C(_0495_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2280_ (.I(_0385_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2281_ (.A1(_0412_),
    .A2(_0476_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2282_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2283_ (.I(_0497_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2284_ (.A1(\ttA_0.data[8][0] ),
    .A2(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2285_ (.A1(_0496_),
    .A2(_0498_),
    .B(_0500_),
    .C(_0495_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2286_ (.I(_0394_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2287_ (.A1(\ttA_0.data[8][1] ),
    .A2(_0499_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2288_ (.A1(_0501_),
    .A2(_0498_),
    .B(_0502_),
    .C(_0495_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2289_ (.I(_0399_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2290_ (.A1(\ttA_0.data[8][2] ),
    .A2(_0499_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2291_ (.A1(_0503_),
    .A2(_0498_),
    .B(_0504_),
    .C(_0495_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2292_ (.I(_0404_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2293_ (.A1(\ttA_0.data[8][3] ),
    .A2(_0499_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2294_ (.I(_0421_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2295_ (.A1(_0505_),
    .A2(_0498_),
    .B(_0506_),
    .C(_0507_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2296_ (.A1(_0379_),
    .A2(_0487_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2297_ (.I(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2298_ (.I(_0508_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2299_ (.A1(\ttA_0.data[5][0] ),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2300_ (.A1(_0496_),
    .A2(_0509_),
    .B(_0511_),
    .C(_0507_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2301_ (.A1(\ttA_0.data[5][1] ),
    .A2(_0510_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2302_ (.A1(_0501_),
    .A2(_0509_),
    .B(_0512_),
    .C(_0507_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2303_ (.A1(\ttA_0.data[5][2] ),
    .A2(_0510_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2304_ (.A1(_0503_),
    .A2(_0509_),
    .B(_0513_),
    .C(_0507_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2305_ (.A1(\ttA_0.data[5][3] ),
    .A2(_0510_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2306_ (.I(_0420_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2307_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2308_ (.A1(_0505_),
    .A2(_0509_),
    .B(_0514_),
    .C(_0516_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2309_ (.A1(_0349_),
    .A2(_0411_),
    .A3(_0375_),
    .A4(_0377_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2310_ (.A1(_0487_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2311_ (.I(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2312_ (.I(_0518_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2313_ (.A1(\ttA_0.data[6][0] ),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2314_ (.A1(_0496_),
    .A2(_0519_),
    .B(_0521_),
    .C(_0516_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2315_ (.A1(\ttA_0.data[6][1] ),
    .A2(_0520_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2316_ (.A1(_0501_),
    .A2(_0519_),
    .B(_0522_),
    .C(_0516_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2317_ (.A1(\ttA_0.data[6][2] ),
    .A2(_0520_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2318_ (.A1(_0503_),
    .A2(_0519_),
    .B(_0523_),
    .C(_0516_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2319_ (.A1(\ttA_0.data[6][3] ),
    .A2(_0520_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2320_ (.I(_0515_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2321_ (.A1(_0505_),
    .A2(_0519_),
    .B(_0524_),
    .C(_0525_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2322_ (.A1(_0412_),
    .A2(_0487_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2323_ (.I(_0526_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2324_ (.I(_0526_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(\ttA_0.data[4][0] ),
    .A2(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2326_ (.A1(_0496_),
    .A2(_0527_),
    .B(_0529_),
    .C(_0525_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2327_ (.A1(\ttA_0.data[4][1] ),
    .A2(_0528_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2328_ (.A1(_0501_),
    .A2(_0527_),
    .B(_0530_),
    .C(_0525_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2329_ (.A1(\ttA_0.data[4][2] ),
    .A2(_0528_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2330_ (.A1(_0503_),
    .A2(_0527_),
    .B(_0531_),
    .C(_0525_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2331_ (.A1(\ttA_0.data[4][3] ),
    .A2(_0528_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2332_ (.I(_0515_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2333_ (.A1(_0505_),
    .A2(_0527_),
    .B(_0532_),
    .C(_0533_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2334_ (.I(_1140_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2335_ (.A1(_1332_),
    .A2(_1396_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2336_ (.I(_0535_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2337_ (.A1(_1104_),
    .A2(_1077_),
    .A3(_1370_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2338_ (.A1(_0256_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2339_ (.A1(_1419_),
    .A2(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2340_ (.A1(_0536_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2341_ (.I(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2342_ (.I(_0540_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2343_ (.A1(\ttA_0.prog[15][0] ),
    .A2(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2344_ (.A1(_0534_),
    .A2(_0541_),
    .B(_0543_),
    .C(_0533_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2345_ (.A1(\ttA_0.prog[15][1] ),
    .A2(_0542_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2346_ (.A1(_0432_),
    .A2(_0541_),
    .B(_0544_),
    .C(_0533_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2347_ (.A1(\ttA_0.prog[15][2] ),
    .A2(_0542_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2348_ (.A1(_0437_),
    .A2(_0541_),
    .B(_0545_),
    .C(_0533_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2349_ (.I(_1180_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2350_ (.A1(\ttA_0.prog[15][3] ),
    .A2(_0542_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2351_ (.I(_0515_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2352_ (.A1(_0546_),
    .A2(_0541_),
    .B(_0547_),
    .C(_0548_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2353_ (.I(_1140_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2354_ (.A1(_1334_),
    .A2(_1396_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2355_ (.A1(_0550_),
    .A2(_0539_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2356_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2357_ (.I(_0551_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2358_ (.I(_1370_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2359_ (.I(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2360_ (.I(_0555_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2361_ (.A1(\ttA_0.prog[14][0] ),
    .A2(_0553_),
    .B(_0000_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2362_ (.A1(_0549_),
    .A2(_0552_),
    .B(_0556_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2363_ (.I(_0555_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2364_ (.A1(\ttA_0.prog[14][1] ),
    .A2(_0553_),
    .B(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2365_ (.A1(_0433_),
    .A2(_0552_),
    .B(_0558_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2366_ (.A1(\ttA_0.prog[14][2] ),
    .A2(_0553_),
    .B(_0557_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2367_ (.A1(_0438_),
    .A2(_0552_),
    .B(_0559_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2368_ (.A1(\ttA_0.prog[14][3] ),
    .A2(_0553_),
    .B(_0557_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2369_ (.A1(_0440_),
    .A2(_0552_),
    .B(_0560_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2370_ (.A1(_1332_),
    .A2(_0376_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2371_ (.A1(_0561_),
    .A2(_0539_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2372_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2373_ (.I(_0562_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2374_ (.A1(\ttA_0.prog[13][0] ),
    .A2(_0564_),
    .B(_0557_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2375_ (.A1(_0549_),
    .A2(_0563_),
    .B(_0565_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2376_ (.I(_0555_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2377_ (.A1(\ttA_0.prog[13][1] ),
    .A2(_0564_),
    .B(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2378_ (.A1(_0433_),
    .A2(_0563_),
    .B(_0567_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2379_ (.A1(\ttA_0.prog[13][2] ),
    .A2(_0564_),
    .B(_0566_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2380_ (.A1(_0438_),
    .A2(_0563_),
    .B(_0568_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2381_ (.A1(\ttA_0.prog[13][3] ),
    .A2(_0564_),
    .B(_0566_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2382_ (.A1(_0440_),
    .A2(_0563_),
    .B(_0569_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2383_ (.A1(_1334_),
    .A2(_0376_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2384_ (.A1(_0570_),
    .A2(_0539_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2385_ (.I(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2386_ (.I(_0571_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2387_ (.A1(\ttA_0.prog[12][0] ),
    .A2(_0573_),
    .B(_0566_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2388_ (.A1(_0549_),
    .A2(_0572_),
    .B(_0574_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2389_ (.I(_0554_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2390_ (.I(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2391_ (.A1(\ttA_0.prog[12][1] ),
    .A2(_0573_),
    .B(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2392_ (.A1(_0423_),
    .A2(_0572_),
    .B(_0577_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2393_ (.A1(\ttA_0.prog[12][2] ),
    .A2(_0573_),
    .B(_0576_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2394_ (.A1(_0428_),
    .A2(_0572_),
    .B(_0578_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2395_ (.A1(\ttA_0.prog[12][3] ),
    .A2(_0573_),
    .B(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2396_ (.A1(_0430_),
    .A2(_0572_),
    .B(_0579_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2397_ (.I(\ttA_0.prog[11][0] ),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2398_ (.I(_0538_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2399_ (.A1(_1420_),
    .A2(_0536_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2400_ (.A1(_0581_),
    .A2(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2401_ (.I(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2402_ (.I(_1176_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2403_ (.I(_0583_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2404_ (.A1(_0585_),
    .A2(_0586_),
    .B(_0576_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2405_ (.A1(_0580_),
    .A2(_0584_),
    .B(_0587_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2406_ (.I(\ttA_0.prog[11][1] ),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2407_ (.I(_0575_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2408_ (.A1(_0452_),
    .A2(_0586_),
    .B(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2409_ (.A1(_0588_),
    .A2(_0584_),
    .B(_0590_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2410_ (.I(\ttA_0.prog[11][2] ),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2411_ (.I(net7),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2412_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2413_ (.A1(_0593_),
    .A2(_0586_),
    .B(_0589_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2414_ (.A1(_0591_),
    .A2(_0584_),
    .B(_0594_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2415_ (.I(\ttA_0.prog[11][3] ),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2416_ (.A1(_1196_),
    .A2(_0586_),
    .B(_0589_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2417_ (.A1(_0595_),
    .A2(_0584_),
    .B(_0596_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2418_ (.I(\ttA_0.prog[10][0] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2419_ (.A1(_1420_),
    .A2(_0550_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2420_ (.A1(_0581_),
    .A2(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2421_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2422_ (.I(_0599_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2423_ (.A1(_0585_),
    .A2(_0601_),
    .B(_0589_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2424_ (.A1(_0597_),
    .A2(_0600_),
    .B(_0602_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2425_ (.I(\ttA_0.prog[10][1] ),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2426_ (.I(_0575_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2427_ (.A1(_0452_),
    .A2(_0601_),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2428_ (.A1(_0603_),
    .A2(_0600_),
    .B(_0605_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2429_ (.I(\ttA_0.prog[10][2] ),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2430_ (.A1(_0593_),
    .A2(_0601_),
    .B(_0604_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2431_ (.A1(_0606_),
    .A2(_0600_),
    .B(_0607_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2432_ (.I(\ttA_0.prog[10][3] ),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2433_ (.A1(_1196_),
    .A2(_0601_),
    .B(_0604_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2434_ (.A1(_0608_),
    .A2(_0600_),
    .B(_0609_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2435_ (.I(\ttA_0.prog[9][0] ),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2436_ (.A1(_1420_),
    .A2(_0561_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2437_ (.A1(_0581_),
    .A2(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2438_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2439_ (.I(_0612_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2440_ (.A1(_0585_),
    .A2(_0614_),
    .B(_0604_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2441_ (.A1(_0610_),
    .A2(_0613_),
    .B(_0615_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2442_ (.I(\ttA_0.prog[9][1] ),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_0575_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2444_ (.A1(_0452_),
    .A2(_0614_),
    .B(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2445_ (.A1(_0616_),
    .A2(_0613_),
    .B(_0618_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2446_ (.I(\ttA_0.prog[9][2] ),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2447_ (.I(net7),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2448_ (.A1(_0620_),
    .A2(_0614_),
    .B(_0617_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2449_ (.A1(_0619_),
    .A2(_0613_),
    .B(_0621_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2450_ (.I(\ttA_0.prog[9][3] ),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2451_ (.I(_1087_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2452_ (.A1(_0623_),
    .A2(_0614_),
    .B(_0617_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2453_ (.A1(_0622_),
    .A2(_0613_),
    .B(_0624_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2454_ (.I(\ttA_0.prog[8][0] ),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2455_ (.A1(_1419_),
    .A2(_0570_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2456_ (.A1(_0581_),
    .A2(_0626_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2457_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2458_ (.I(_0627_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2459_ (.A1(_0585_),
    .A2(_0629_),
    .B(_0617_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2460_ (.A1(_0625_),
    .A2(_0628_),
    .B(_0630_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2461_ (.I(\ttA_0.prog[8][1] ),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2462_ (.I(_1123_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2463_ (.I(_0554_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2464_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2465_ (.A1(_0632_),
    .A2(_0629_),
    .B(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2466_ (.A1(_0631_),
    .A2(_0628_),
    .B(_0635_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2467_ (.I(\ttA_0.prog[8][2] ),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2468_ (.A1(_0620_),
    .A2(_0629_),
    .B(_0634_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2469_ (.A1(_0636_),
    .A2(_0628_),
    .B(_0637_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2470_ (.I(\ttA_0.prog[8][3] ),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2471_ (.A1(_0623_),
    .A2(_0629_),
    .B(_0634_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2472_ (.A1(_0638_),
    .A2(_0628_),
    .B(_0639_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2473_ (.I(\ttA_0.prog[7][0] ),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2474_ (.A1(_0318_),
    .A2(_0535_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2475_ (.I(_0537_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2476_ (.A1(_1434_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2477_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2478_ (.A1(_0641_),
    .A2(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2479_ (.I(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2480_ (.I(_1176_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2481_ (.I(_0645_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2482_ (.A1(_0647_),
    .A2(_0648_),
    .B(_0634_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2483_ (.A1(_0640_),
    .A2(_0646_),
    .B(_0649_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2484_ (.I(\ttA_0.prog[7][1] ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2485_ (.I(_0633_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2486_ (.A1(_0632_),
    .A2(_0648_),
    .B(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2487_ (.A1(_0650_),
    .A2(_0646_),
    .B(_0652_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2488_ (.I(\ttA_0.prog[7][2] ),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0620_),
    .A2(_0648_),
    .B(_0651_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2490_ (.A1(_0653_),
    .A2(_0646_),
    .B(_0654_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2491_ (.I(\ttA_0.prog[7][3] ),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2492_ (.A1(_0623_),
    .A2(_0648_),
    .B(_0651_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2493_ (.A1(_0655_),
    .A2(_0646_),
    .B(_0656_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(_1419_),
    .A2(_0256_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2495_ (.A1(_0550_),
    .A2(_0657_),
    .A3(_0642_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2496_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2497_ (.I(_0658_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2498_ (.A1(\ttA_0.prog[6][0] ),
    .A2(_0660_),
    .B(_0651_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2499_ (.A1(_0534_),
    .A2(_0659_),
    .B(_0661_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2500_ (.I(_0633_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2501_ (.A1(\ttA_0.prog[6][1] ),
    .A2(_0660_),
    .B(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2502_ (.A1(_0423_),
    .A2(_0659_),
    .B(_0663_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2503_ (.A1(\ttA_0.prog[6][2] ),
    .A2(_0660_),
    .B(_0662_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2504_ (.A1(_0428_),
    .A2(_0659_),
    .B(_0664_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2505_ (.A1(\ttA_0.prog[6][3] ),
    .A2(_0660_),
    .B(_0662_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2506_ (.A1(_0430_),
    .A2(_0659_),
    .B(_0665_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2507_ (.A1(_0561_),
    .A2(_0657_),
    .A3(_0642_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2508_ (.I(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2509_ (.I(_0666_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2510_ (.A1(\ttA_0.prog[5][0] ),
    .A2(_0668_),
    .B(_0662_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2511_ (.A1(_0534_),
    .A2(_0667_),
    .B(_0669_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2512_ (.I(_0633_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2513_ (.A1(\ttA_0.prog[5][1] ),
    .A2(_0668_),
    .B(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2514_ (.A1(_0423_),
    .A2(_0667_),
    .B(_0671_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2515_ (.A1(\ttA_0.prog[5][2] ),
    .A2(_0668_),
    .B(_0670_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2516_ (.A1(_0428_),
    .A2(_0667_),
    .B(_0672_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2517_ (.A1(\ttA_0.prog[5][3] ),
    .A2(_0668_),
    .B(_0670_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2518_ (.A1(_0430_),
    .A2(_0667_),
    .B(_0673_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2519_ (.A1(_0570_),
    .A2(_0657_),
    .A3(_0642_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2520_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2521_ (.I(_0674_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2522_ (.A1(\ttA_0.prog[4][0] ),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2523_ (.A1(_0534_),
    .A2(_0675_),
    .B(_0677_),
    .C(_0548_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2524_ (.A1(\ttA_0.prog[4][1] ),
    .A2(_0676_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2525_ (.A1(_0432_),
    .A2(_0675_),
    .B(_0678_),
    .C(_0548_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2526_ (.A1(\ttA_0.prog[4][2] ),
    .A2(_0676_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2527_ (.A1(_0437_),
    .A2(_0675_),
    .B(_0679_),
    .C(_0548_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2528_ (.A1(\ttA_0.prog[4][3] ),
    .A2(_0676_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2529_ (.I(_0420_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2530_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2531_ (.A1(_0546_),
    .A2(_0675_),
    .B(_0680_),
    .C(_0682_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2532_ (.I(_1223_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2533_ (.A1(\ttA_1.top.data[7][0] ),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2534_ (.A1(_0432_),
    .A2(_0683_),
    .B(_0684_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2535_ (.A1(\ttA_1.top.data[7][1] ),
    .A2(_1223_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2536_ (.A1(_0437_),
    .A2(_0683_),
    .B(_0685_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2537_ (.A1(\ttA_1.top.data[7][2] ),
    .A2(_1223_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2538_ (.A1(_0546_),
    .A2(_0683_),
    .B(_0686_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2539_ (.I(\ttA_0.io_out[4] ),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2540_ (.I(_0687_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2541_ (.A1(_0273_),
    .A2(_0283_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2542_ (.I(_0311_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2543_ (.A1(_1433_),
    .A2(_0296_),
    .A3(_0301_),
    .B1(_0286_),
    .B2(_0290_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2544_ (.I(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2545_ (.A1(_0690_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2546_ (.A1(_0689_),
    .A2(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2547_ (.A1(_0689_),
    .A2(_0690_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2548_ (.I(_0273_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2549_ (.A1(_0280_),
    .A2(_0282_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2550_ (.A1(_1432_),
    .A2(_0276_),
    .A3(_0278_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2551_ (.A1(_0696_),
    .A2(_0697_),
    .A3(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2552_ (.A1(_0693_),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2553_ (.A1(_0695_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2554_ (.A1(_0291_),
    .A2(_0302_),
    .B(_0694_),
    .C(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2555_ (.A1(_1402_),
    .A2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2556_ (.I(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2557_ (.I(_0362_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2558_ (.A1(_0695_),
    .A2(_0700_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2559_ (.A1(_0705_),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2560_ (.A1(_1476_),
    .A2(_0374_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2561_ (.A1(\ttA_0.io_out[7] ),
    .A2(_0326_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2562_ (.A1(_1500_),
    .A2(_0343_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2563_ (.A1(_1470_),
    .A2(_0359_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2564_ (.A1(_0708_),
    .A2(_0709_),
    .A3(_0710_),
    .A4(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2565_ (.A1(_0693_),
    .A2(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2566_ (.I(_0312_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2567_ (.A1(_1508_),
    .A2(_1501_),
    .A3(_0391_),
    .A4(_1470_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2568_ (.A1(_0326_),
    .A2(_0473_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2569_ (.A1(_0359_),
    .A2(_0373_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2570_ (.A1(_0715_),
    .A2(_0716_),
    .A3(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2571_ (.I(_0690_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2572_ (.A1(_0719_),
    .A2(_0692_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2573_ (.A1(_0690_),
    .A2(_0692_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2574_ (.A1(_0716_),
    .A2(_0717_),
    .B(_0721_),
    .C(_0715_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2575_ (.A1(_0714_),
    .A2(_0718_),
    .B1(_0712_),
    .B2(_0720_),
    .C(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2576_ (.A1(_0697_),
    .A2(_0698_),
    .B1(_0713_),
    .B2(_0723_),
    .C(_0696_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2577_ (.A1(_0696_),
    .A2(_0283_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2578_ (.A1(_0687_),
    .A2(_0362_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2579_ (.A1(_0720_),
    .A2(_0715_),
    .B1(_0726_),
    .B2(_0714_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2580_ (.A1(_0693_),
    .A2(_0725_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2581_ (.A1(_0688_),
    .A2(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2582_ (.A1(_0725_),
    .A2(_0727_),
    .B(_0729_),
    .C(_0701_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2583_ (.A1(_0326_),
    .A2(_0473_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2584_ (.I(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2585_ (.I(_0374_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2586_ (.I(\ttA_0.io_out[6] ),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2587_ (.I(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2588_ (.I(_0409_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2589_ (.A1(_1508_),
    .A2(_0409_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2590_ (.A1(_0735_),
    .A2(_0736_),
    .B(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2591_ (.A1(_1471_),
    .A2(_0362_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2592_ (.A1(_0391_),
    .A2(_0409_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2593_ (.I(_0325_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2594_ (.A1(_0739_),
    .A2(_0740_),
    .B(_0741_),
    .C(_0733_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2595_ (.A1(_0733_),
    .A2(_0738_),
    .B(_0742_),
    .C(_0731_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2596_ (.A1(_0273_),
    .A2(_0697_),
    .A3(_0698_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2597_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2598_ (.A1(_0745_),
    .A2(_0720_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2599_ (.A1(_1509_),
    .A2(_0732_),
    .B(_0743_),
    .C(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2600_ (.I(_0741_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2601_ (.A1(_0748_),
    .A2(_0739_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2602_ (.I(_0373_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2603_ (.I(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2604_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2605_ (.A1(_0714_),
    .A2(_0745_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2606_ (.A1(_0753_),
    .A2(_0731_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2607_ (.A1(_0752_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2608_ (.I(_0694_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2609_ (.A1(_0721_),
    .A2(_0725_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2610_ (.A1(_0687_),
    .A2(_0361_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2611_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2612_ (.A1(_0311_),
    .A2(_0691_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2613_ (.A1(_0745_),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2614_ (.A1(_0689_),
    .A2(_0719_),
    .A3(_0692_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2615_ (.A1(_0762_),
    .A2(_0711_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2616_ (.A1(_0749_),
    .A2(_0755_),
    .B(_0759_),
    .C(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2617_ (.A1(_0724_),
    .A2(_0730_),
    .A3(_0747_),
    .A4(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2618_ (.A1(_0707_),
    .A2(_0765_),
    .B(_0704_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2619_ (.A1(_0688_),
    .A2(_0704_),
    .B(_0766_),
    .C(_0682_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2620_ (.I(_0703_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2621_ (.A1(_1470_),
    .A2(_0361_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2622_ (.A1(_0745_),
    .A2(_0760_),
    .B(_0360_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2623_ (.A1(_1477_),
    .A2(_0750_),
    .A3(_0769_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2624_ (.A1(_0768_),
    .A2(_0770_),
    .B(_0762_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2625_ (.A1(_0768_),
    .A2(_0770_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2626_ (.A1(_0392_),
    .A2(_0705_),
    .B(_0758_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2627_ (.A1(_0688_),
    .A2(_0752_),
    .B(_0740_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2628_ (.A1(\ttA_0.io_out[5] ),
    .A2(_0373_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2629_ (.A1(_0775_),
    .A2(_0758_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2630_ (.A1(_0756_),
    .A2(_0774_),
    .A3(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2631_ (.I(_0733_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2632_ (.A1(_0696_),
    .A2(_0283_),
    .A3(_0714_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2633_ (.A1(_0391_),
    .A2(_0778_),
    .B(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(_0701_),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2635_ (.A1(_0775_),
    .A2(_0757_),
    .B1(_0728_),
    .B2(_1477_),
    .C(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2636_ (.A1(_0755_),
    .A2(_0773_),
    .B(_0777_),
    .C(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2637_ (.I(_0733_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2638_ (.A1(_0402_),
    .A2(_0705_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2639_ (.I(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2640_ (.A1(_0392_),
    .A2(_0705_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2641_ (.A1(_1502_),
    .A2(_0736_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2642_ (.A1(_0787_),
    .A2(_0788_),
    .B(_0748_),
    .C(_0778_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2643_ (.A1(_0784_),
    .A2(_0786_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2644_ (.A1(_0746_),
    .A2(_0732_),
    .A3(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2645_ (.A1(_0772_),
    .A2(_0783_),
    .A3(_0791_),
    .B1(_0701_),
    .B2(_0784_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2646_ (.A1(_0392_),
    .A2(_0767_),
    .B(_0670_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2647_ (.A1(_0767_),
    .A2(_0792_),
    .B(_0793_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2648_ (.A1(_0751_),
    .A2(_0769_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_0751_),
    .A2(_0769_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2650_ (.A1(_1477_),
    .A2(_0794_),
    .A3(_0795_),
    .B1(_0770_),
    .B2(_0768_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2651_ (.A1(_0744_),
    .A2(_0760_),
    .B(_0717_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2652_ (.A1(_0344_),
    .A2(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2653_ (.A1(_1500_),
    .A2(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2654_ (.A1(_0699_),
    .A2(_0721_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2655_ (.A1(_0284_),
    .A2(_0720_),
    .B(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2656_ (.A1(_0796_),
    .A2(_0799_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2657_ (.A1(_0796_),
    .A2(_0799_),
    .B(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2658_ (.A1(_0734_),
    .A2(_0361_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(\ttA_0.io_out[4] ),
    .A2(_0342_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2660_ (.A1(_0775_),
    .A2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2661_ (.A1(_0804_),
    .A2(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2662_ (.A1(_0776_),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2663_ (.I(_0473_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2664_ (.A1(_0778_),
    .A2(_0746_),
    .A3(_0732_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2665_ (.A1(_0735_),
    .A2(_0728_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2666_ (.A1(_1502_),
    .A2(_0809_),
    .A3(_0757_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2667_ (.A1(_1501_),
    .A2(_0809_),
    .B(_0779_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2668_ (.A1(_0811_),
    .A2(_0812_),
    .A3(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2669_ (.A1(_0809_),
    .A2(_0706_),
    .B1(_0738_),
    .B2(_0810_),
    .C(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2670_ (.I(_0741_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2671_ (.A1(_0816_),
    .A2(_0740_),
    .B(_0752_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2672_ (.A1(_0735_),
    .A2(_0816_),
    .A3(_0736_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_0778_),
    .A2(_0749_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2674_ (.A1(_0817_),
    .A2(_0818_),
    .B(_0819_),
    .C(_0754_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2675_ (.A1(_0767_),
    .A2(_0815_),
    .A3(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2676_ (.A1(_0756_),
    .A2(_0808_),
    .B(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2677_ (.I(_0389_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2678_ (.A1(_0735_),
    .A2(_0704_),
    .B1(_0803_),
    .B2(_0822_),
    .C(_0823_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2679_ (.A1(_1501_),
    .A2(_0798_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2680_ (.A1(_0796_),
    .A2(_0799_),
    .B(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2681_ (.A1(_0344_),
    .A2(_0717_),
    .B(_0800_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2682_ (.A1(_0709_),
    .A2(_0825_),
    .A3(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2683_ (.A1(_0801_),
    .A2(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2684_ (.A1(_0775_),
    .A2(_0758_),
    .A3(_0807_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(_1471_),
    .A2(_0741_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2686_ (.A1(_0804_),
    .A2(_0806_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2687_ (.A1(_0687_),
    .A2(_0751_),
    .B(_0343_),
    .C(_1476_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_1500_),
    .A2(_0374_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2689_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2690_ (.A1(_0830_),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2691_ (.A1(_0737_),
    .A2(_0829_),
    .A3(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2692_ (.A1(_0402_),
    .A2(_0748_),
    .A3(_0757_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2693_ (.A1(_0402_),
    .A2(_0748_),
    .B(_0779_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2694_ (.A1(_1509_),
    .A2(_0728_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2695_ (.A1(_0837_),
    .A2(_0838_),
    .A3(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2696_ (.A1(_0816_),
    .A2(_0706_),
    .B1(_0786_),
    .B2(_0810_),
    .C(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2697_ (.A1(_0784_),
    .A2(_0716_),
    .A3(_0773_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2698_ (.A1(_0752_),
    .A2(_0716_),
    .A3(_0785_),
    .A4(_0788_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2699_ (.A1(_0688_),
    .A2(_0732_),
    .B(_0753_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2700_ (.A1(_0842_),
    .A2(_0843_),
    .A3(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2701_ (.A1(_0767_),
    .A2(_0841_),
    .A3(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2702_ (.A1(_0756_),
    .A2(_0836_),
    .B(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2703_ (.I(_1377_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2704_ (.A1(_1509_),
    .A2(_0704_),
    .B1(_0828_),
    .B2(_0847_),
    .C(_0848_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2705_ (.I(_0385_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2706_ (.A1(_0328_),
    .A2(_0347_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2707_ (.A1(_0517_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2708_ (.I(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2709_ (.I(_0851_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2710_ (.A1(\ttA_0.data[14][0] ),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2711_ (.A1(_0849_),
    .A2(_0852_),
    .B(_0854_),
    .C(_0682_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2712_ (.I(_0394_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2713_ (.A1(\ttA_0.data[14][1] ),
    .A2(_0853_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2714_ (.A1(_0855_),
    .A2(_0852_),
    .B(_0856_),
    .C(_0682_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2715_ (.I(_0399_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2716_ (.A1(\ttA_0.data[14][2] ),
    .A2(_0853_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2717_ (.I(_0681_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2718_ (.A1(_0857_),
    .A2(_0852_),
    .B(_0858_),
    .C(_0859_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2719_ (.I(_0404_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(\ttA_0.data[14][3] ),
    .A2(_0853_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2721_ (.A1(_0860_),
    .A2(_0852_),
    .B(_0861_),
    .C(_0859_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2722_ (.I(_0848_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2723_ (.I(_0862_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2724_ (.I(_0862_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2725_ (.A1(_0348_),
    .A2(_0485_),
    .A3(_0486_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2726_ (.I(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2727_ (.I(_0863_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2728_ (.A1(\ttA_0.data[3][0] ),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2729_ (.A1(_0849_),
    .A2(_0864_),
    .B(_0866_),
    .C(_0859_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2730_ (.A1(\ttA_0.data[3][1] ),
    .A2(_0865_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2731_ (.A1(_0855_),
    .A2(_0864_),
    .B(_0867_),
    .C(_0859_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2732_ (.A1(\ttA_0.data[3][2] ),
    .A2(_0865_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_0681_),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2734_ (.A1(_0857_),
    .A2(_0864_),
    .B(_0868_),
    .C(_0869_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2735_ (.A1(\ttA_0.data[3][3] ),
    .A2(_0865_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2736_ (.A1(_0860_),
    .A2(_0864_),
    .B(_0870_),
    .C(_0869_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2737_ (.A1(_0412_),
    .A2(_0850_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2738_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2739_ (.I(_0871_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2740_ (.A1(\ttA_0.data[12][0] ),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2741_ (.A1(_0849_),
    .A2(_0872_),
    .B(_0874_),
    .C(_0869_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2742_ (.A1(\ttA_0.data[12][1] ),
    .A2(_0873_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2743_ (.A1(_0855_),
    .A2(_0872_),
    .B(_0875_),
    .C(_0869_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2744_ (.A1(\ttA_0.data[12][2] ),
    .A2(_0873_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2745_ (.I(_0681_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2746_ (.A1(_0857_),
    .A2(_0872_),
    .B(_0876_),
    .C(_0877_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2747_ (.A1(\ttA_0.data[12][3] ),
    .A2(_0873_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2748_ (.A1(_0860_),
    .A2(_0872_),
    .B(_0878_),
    .C(_0877_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2749_ (.A1(_0485_),
    .A2(_0486_),
    .A3(_0850_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2750_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2751_ (.I(_0879_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2752_ (.A1(\ttA_0.data[15][0] ),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2753_ (.A1(_0849_),
    .A2(_0880_),
    .B(_0882_),
    .C(_0877_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2754_ (.A1(\ttA_0.data[15][1] ),
    .A2(_0881_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2755_ (.A1(_0855_),
    .A2(_0880_),
    .B(_0883_),
    .C(_0877_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2756_ (.A1(\ttA_0.data[15][2] ),
    .A2(_0881_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2757_ (.I(_0420_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2758_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2759_ (.A1(_0857_),
    .A2(_0880_),
    .B(_0884_),
    .C(_0886_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2760_ (.A1(\ttA_0.data[15][3] ),
    .A2(_0881_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2761_ (.A1(_0860_),
    .A2(_0880_),
    .B(_0887_),
    .C(_0886_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2762_ (.I(_0385_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_0476_),
    .A2(_0517_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2764_ (.I(_0889_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2765_ (.I(_0889_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2766_ (.A1(\ttA_0.data[10][0] ),
    .A2(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2767_ (.A1(_0888_),
    .A2(_0890_),
    .B(_0892_),
    .C(_0886_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2768_ (.I(_0394_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2769_ (.A1(\ttA_0.data[10][1] ),
    .A2(_0891_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2770_ (.A1(_0893_),
    .A2(_0890_),
    .B(_0894_),
    .C(_0886_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2771_ (.I(_0399_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(\ttA_0.data[10][2] ),
    .A2(_0891_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2773_ (.I(_0885_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2774_ (.A1(_0895_),
    .A2(_0890_),
    .B(_0896_),
    .C(_0897_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2775_ (.I(_0404_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2776_ (.A1(\ttA_0.data[10][3] ),
    .A2(_0891_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2777_ (.A1(_0898_),
    .A2(_0890_),
    .B(_0899_),
    .C(_0897_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2778_ (.I(\ttA_0.prog[3][0] ),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2779_ (.A1(_0582_),
    .A2(_0644_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2780_ (.I(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2781_ (.I(_0901_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2782_ (.I(_0554_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2783_ (.I(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2784_ (.A1(_0647_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2785_ (.A1(_0900_),
    .A2(_0902_),
    .B(_0906_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2786_ (.I(\ttA_0.prog[3][1] ),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2787_ (.A1(_0632_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2788_ (.A1(_0907_),
    .A2(_0902_),
    .B(_0908_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2789_ (.I(\ttA_0.prog[3][2] ),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2790_ (.A1(_0620_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2791_ (.A1(_0909_),
    .A2(_0902_),
    .B(_0910_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2792_ (.I(\ttA_0.prog[3][3] ),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2793_ (.A1(_0623_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2794_ (.A1(_0911_),
    .A2(_0902_),
    .B(_0912_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2795_ (.I(_1368_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2796_ (.I(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2797_ (.I(_0914_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2798_ (.I(_0914_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2799_ (.I(_0914_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2800_ (.I(_0914_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2801_ (.I(_1368_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2802_ (.I(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2803_ (.I(_0916_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2804_ (.I(_0916_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2805_ (.I(_0916_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2806_ (.I(_0916_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2807_ (.I(_0915_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2808_ (.I(_0917_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2809_ (.I(_0917_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2810_ (.I(_0917_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2811_ (.A1(_0348_),
    .A2(_0517_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2812_ (.I(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2813_ (.I(_0918_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2814_ (.A1(\ttA_0.data[2][0] ),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2815_ (.A1(_0888_),
    .A2(_0919_),
    .B(_0921_),
    .C(_0897_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(\ttA_0.data[2][1] ),
    .A2(_0920_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2817_ (.A1(_0893_),
    .A2(_0919_),
    .B(_0922_),
    .C(_0897_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2818_ (.A1(\ttA_0.data[2][2] ),
    .A2(_0920_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2819_ (.I(_0885_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2820_ (.A1(_0895_),
    .A2(_0919_),
    .B(_0923_),
    .C(_0924_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2821_ (.A1(\ttA_0.data[2][3] ),
    .A2(_0920_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2822_ (.A1(_0898_),
    .A2(_0919_),
    .B(_0925_),
    .C(_0924_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2823_ (.I(_0917_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2824_ (.I(_0915_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2825_ (.I(_0926_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2826_ (.I(_0926_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2827_ (.I(_0926_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2828_ (.I(_0926_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2829_ (.I(_0915_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2830_ (.I(_0927_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2831_ (.I(_0927_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2832_ (.I(_0927_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2833_ (.I(_0407_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2834_ (.A1(_0440_),
    .A2(_0928_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2835_ (.I(_0862_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2836_ (.I(\ttA_4.counter[4] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2837_ (.I(\ttA_4.counter[3] ),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2838_ (.I(\ttA_4.active_duty[3] ),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2839_ (.I(\ttA_4.active_duty[2] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2840_ (.I(\ttA_4.counter[1] ),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2841_ (.I(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2842_ (.I(\ttA_4.counter[0] ),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2843_ (.A1(\ttA_4.active_duty[1] ),
    .A2(_0934_),
    .B(\ttA_4.active_duty[0] ),
    .C(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2844_ (.I(\ttA_4.counter[2] ),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2845_ (.A1(\ttA_4.active_duty[2] ),
    .A2(_0937_),
    .B1(\ttA_4.active_duty[1] ),
    .B2(_0934_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2846_ (.A1(_0931_),
    .A2(\ttA_4.counter[3] ),
    .B1(_0932_),
    .B2(\ttA_4.counter[2] ),
    .C1(_0936_),
    .C2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2847_ (.A1(\ttA_4.active_duty[4] ),
    .A2(_0929_),
    .B1(\ttA_4.active_duty[3] ),
    .B2(_0930_),
    .C(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2848_ (.I(\ttA_4.active_duty[5] ),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2849_ (.I(\ttA_4.active_duty[4] ),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2850_ (.A1(_0941_),
    .A2(\ttA_4.counter[5] ),
    .B1(_0942_),
    .B2(\ttA_4.counter[4] ),
    .C(_0389_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2851_ (.I(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(\ttA_4.active_duty[5] ),
    .A2(_0555_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2853_ (.A1(_0407_),
    .A2(\ttA_4.pwm_signal ),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2854_ (.A1(_0940_),
    .A2(_0944_),
    .B1(_0945_),
    .B2(\ttA_4.counter[5] ),
    .C(_0946_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2855_ (.I(\ttA_0.prog[2][0] ),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2856_ (.A1(_0598_),
    .A2(_0644_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2857_ (.I(_0948_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2858_ (.I(_0948_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2859_ (.I(_0904_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2860_ (.A1(_0647_),
    .A2(_0950_),
    .B(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2861_ (.A1(_0947_),
    .A2(_0949_),
    .B(_0952_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2862_ (.I(\ttA_0.prog[2][1] ),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2863_ (.A1(_0632_),
    .A2(_0950_),
    .B(_0951_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2864_ (.A1(_0953_),
    .A2(_0949_),
    .B(_0954_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2865_ (.I(\ttA_0.prog[2][2] ),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2866_ (.A1(_0592_),
    .A2(_0950_),
    .B(_0951_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2867_ (.A1(_0955_),
    .A2(_0949_),
    .B(_0956_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2868_ (.I(\ttA_0.prog[2][3] ),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_1088_),
    .A2(_0950_),
    .B(_0951_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2870_ (.A1(_0957_),
    .A2(_0949_),
    .B(_0958_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2871_ (.I(_0927_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2872_ (.I(_0913_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2873_ (.I(_0913_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2874_ (.I(_0913_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2875_ (.A1(_1401_),
    .A2(_1345_),
    .A3(_1355_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2876_ (.I(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2877_ (.A1(_0003_),
    .A2(_1422_),
    .B(_0960_),
    .C(_1386_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2878_ (.A1(net12),
    .A2(_1288_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2879_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2880_ (.A1(net13),
    .A2(_1281_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2881_ (.A1(\beepboop.inst.counter[0] ),
    .A2(_0962_),
    .A3(_0963_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2882_ (.I(\ttA_0.prog[1][0] ),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2883_ (.A1(_0611_),
    .A2(_0644_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2884_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2885_ (.I(_0965_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2886_ (.I(_0904_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2887_ (.A1(_0647_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2888_ (.A1(_0964_),
    .A2(_0966_),
    .B(_0969_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2889_ (.I(\ttA_0.prog[1][1] ),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2890_ (.A1(_1205_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2891_ (.A1(_0970_),
    .A2(_0966_),
    .B(_0971_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2892_ (.I(\ttA_0.prog[1][2] ),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2893_ (.A1(_0592_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2894_ (.A1(_0972_),
    .A2(_0966_),
    .B(_0973_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2895_ (.I(\ttA_0.prog[1][3] ),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2896_ (.A1(_1088_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2897_ (.A1(_0974_),
    .A2(_0966_),
    .B(_0975_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2898_ (.I(\ttA_0.prog[0][0] ),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2899_ (.A1(_0626_),
    .A2(_0643_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2900_ (.I(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2901_ (.I(_0977_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2902_ (.I(_0904_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2903_ (.A1(_1198_),
    .A2(_0979_),
    .B(_0980_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2904_ (.A1(_0976_),
    .A2(_0978_),
    .B(_0981_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2905_ (.I(\ttA_0.prog[0][1] ),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2906_ (.A1(_1205_),
    .A2(_0979_),
    .B(_0980_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2907_ (.A1(_0982_),
    .A2(_0978_),
    .B(_0983_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2908_ (.I(\ttA_0.prog[0][2] ),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2909_ (.A1(_0592_),
    .A2(_0979_),
    .B(_0980_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2910_ (.A1(_0984_),
    .A2(_0978_),
    .B(_0985_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2911_ (.I(\ttA_0.prog[0][3] ),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2912_ (.A1(_1088_),
    .A2(_0979_),
    .B(_0980_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2913_ (.A1(_0986_),
    .A2(_0978_),
    .B(_0987_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2914_ (.I(\ttA_4.counter[0] ),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2915_ (.A1(_0988_),
    .A2(_0928_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2916_ (.A1(\ttA_4.counter[5] ),
    .A2(\ttA_4.counter[4] ),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2917_ (.A1(_0930_),
    .A2(_0937_),
    .A3(_0934_),
    .A4(_0988_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2918_ (.A1(_0989_),
    .A2(_0990_),
    .B(_1401_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2919_ (.I(_0991_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2920_ (.A1(_0934_),
    .A2(_0988_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2921_ (.A1(_0992_),
    .A2(_0993_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2922_ (.A1(_0937_),
    .A2(_0933_),
    .A3(_0935_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2923_ (.A1(\ttA_4.counter[1] ),
    .A2(_0988_),
    .B(\ttA_4.counter[2] ),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2924_ (.A1(_0992_),
    .A2(_0994_),
    .A3(_0995_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2925_ (.A1(\ttA_4.counter[3] ),
    .A2(_0994_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2926_ (.A1(\ttA_4.counter[3] ),
    .A2(_0994_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2927_ (.A1(_0991_),
    .A2(_0996_),
    .A3(_0997_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2928_ (.A1(_0929_),
    .A2(_0996_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2929_ (.A1(_0992_),
    .A2(_0998_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2930_ (.A1(\ttA_4.counter[4] ),
    .A2(_0996_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2931_ (.A1(\ttA_4.counter[5] ),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2932_ (.A1(_0992_),
    .A2(_1000_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2933_ (.A1(_0379_),
    .A2(_0850_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2934_ (.I(_1001_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2935_ (.I(_1001_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2936_ (.A1(\ttA_0.data[13][0] ),
    .A2(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2937_ (.A1(_0888_),
    .A2(_1002_),
    .B(_1004_),
    .C(_0924_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2938_ (.A1(\ttA_0.data[13][1] ),
    .A2(_1003_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2939_ (.A1(_0893_),
    .A2(_1002_),
    .B(_1005_),
    .C(_0924_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2940_ (.A1(\ttA_0.data[13][2] ),
    .A2(_1003_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2941_ (.I(_0885_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2942_ (.A1(_0895_),
    .A2(_1002_),
    .B(_1006_),
    .C(_1007_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2943_ (.A1(\ttA_0.data[13][3] ),
    .A2(_1003_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2944_ (.A1(_0898_),
    .A2(_1002_),
    .B(_1008_),
    .C(_1007_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2945_ (.A1(_1266_),
    .A2(_1256_),
    .B(_0389_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2946_ (.A1(\ttA_4.active_duty[0] ),
    .A2(_0000_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2947_ (.A1(_0003_),
    .A2(_1009_),
    .B(_1010_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2948_ (.A1(\ttA_4.active_duty[1] ),
    .A2(_0823_),
    .B1(_1009_),
    .B2(_1425_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2949_ (.I(_1011_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2950_ (.I(_0407_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2951_ (.A1(_0932_),
    .A2(_1012_),
    .B1(_1009_),
    .B2(_0549_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2952_ (.A1(_0931_),
    .A2(_0390_),
    .B1(_1009_),
    .B2(_0433_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2953_ (.A1(_0593_),
    .A2(_0848_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2954_ (.A1(_0942_),
    .A2(_0928_),
    .B(_1013_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2955_ (.A1(_0546_),
    .A2(_0000_),
    .B(_0945_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2956_ (.I(_1376_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2957_ (.A1(\ttA_0.lastdata3 ),
    .A2(_0700_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2958_ (.A1(_1402_),
    .A2(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2959_ (.A1(_1368_),
    .A2(_1015_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2960_ (.A1(_1425_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2961_ (.A1(_1198_),
    .A2(_1014_),
    .B1(_0736_),
    .B2(_1016_),
    .C1(_1018_),
    .C2(_1334_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2962_ (.A1(_1012_),
    .A2(_1019_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2963_ (.A1(_0570_),
    .A2(_0536_),
    .A3(_1018_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2964_ (.A1(_1205_),
    .A2(_1014_),
    .B1(_0784_),
    .B2(_1016_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2965_ (.A1(_1020_),
    .A2(_1021_),
    .B(_0928_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2966_ (.A1(_0593_),
    .A2(_1014_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2967_ (.A1(_0318_),
    .A2(_0536_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2968_ (.A1(_0809_),
    .A2(_1016_),
    .B1(_1023_),
    .B2(_1018_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2969_ (.A1(_1022_),
    .A2(_1024_),
    .B(_1012_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2970_ (.A1(_1434_),
    .A2(_0641_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2971_ (.A1(_1122_),
    .A2(_1014_),
    .B1(_0816_),
    .B2(_1016_),
    .C1(_1025_),
    .C2(_1018_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2972_ (.A1(_1012_),
    .A2(_1026_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2973_ (.A1(_0485_),
    .A2(_0486_),
    .A3(_0476_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2974_ (.I(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2975_ (.I(_1027_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2976_ (.A1(\ttA_0.data[11][0] ),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2977_ (.A1(_0888_),
    .A2(_1028_),
    .B(_1030_),
    .C(_1007_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2978_ (.A1(\ttA_0.data[11][1] ),
    .A2(_1029_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2979_ (.A1(_0893_),
    .A2(_1028_),
    .B(_1031_),
    .C(_1007_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2980_ (.A1(\ttA_0.data[11][2] ),
    .A2(_1029_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2981_ (.A1(_0895_),
    .A2(_1028_),
    .B(_1032_),
    .C(_0823_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2982_ (.A1(\ttA_0.data[11][3] ),
    .A2(_1029_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2983_ (.A1(_0898_),
    .A2(_1028_),
    .B(_1033_),
    .C(_0823_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2984_ (.A1(\ttA_6.counter[1] ),
    .A2(_1386_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2985_ (.I(_0959_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2986_ (.A1(\ttA_6.counter[1] ),
    .A2(\ttA_6.counter[0] ),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2987_ (.I(_1036_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2988_ (.A1(_1034_),
    .A2(_1035_),
    .A3(_1037_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2989_ (.A1(_1385_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2990_ (.A1(_1035_),
    .A2(_1038_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2991_ (.I(_0959_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2992_ (.A1(_1438_),
    .A2(_1037_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2993_ (.A1(_1385_),
    .A2(_1037_),
    .B(_1358_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2994_ (.A1(_1039_),
    .A2(_1040_),
    .A3(_1041_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2995_ (.A1(\ttA_6.counter[4] ),
    .A2(_1437_),
    .A3(_1036_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2996_ (.A1(_1448_),
    .A2(_1040_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2997_ (.A1(_1039_),
    .A2(_1042_),
    .A3(_1043_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2998_ (.A1(\ttA_6.counter[5] ),
    .A2(_1042_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2999_ (.A1(_1447_),
    .A2(_1042_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3000_ (.A1(_1039_),
    .A2(_1044_),
    .A3(_1045_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3001_ (.A1(\ttA_6.counter[6] ),
    .A2(_1044_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3002_ (.A1(_1456_),
    .A2(_1044_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3003_ (.A1(_1039_),
    .A2(_1046_),
    .A3(_1047_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3004_ (.A1(_1387_),
    .A2(_1046_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3005_ (.A1(\ttA_6.counter[7] ),
    .A2(_1046_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3006_ (.A1(_0960_),
    .A2(_1048_),
    .A3(_1049_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3007_ (.A1(_1436_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3008_ (.A1(\ttA_6.counter[8] ),
    .A2(_1049_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3009_ (.A1(_0960_),
    .A2(_1050_),
    .A3(_1051_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3010_ (.A1(_1441_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3011_ (.A1(_1441_),
    .A2(_1051_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3012_ (.A1(_0960_),
    .A2(_1052_),
    .A3(_1053_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3013_ (.A1(_1435_),
    .A2(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3014_ (.A1(_1035_),
    .A2(_1054_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3015_ (.A1(\ttA_6.counter[10] ),
    .A2(_1053_),
    .B(_1346_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3016_ (.A1(_1035_),
    .A2(_1055_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3017_ (.I(_0862_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3018_ (.I(_0848_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3019_ (.I(_1056_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3020_ (.I(_1056_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3021_ (.I(_1056_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3022_ (.I(_1056_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3023_ (.A1(\beepboop.inst.counter[1] ),
    .A2(\beepboop.inst.counter[0] ),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3024_ (.A1(_1279_),
    .A2(_0962_),
    .A3(_1057_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3025_ (.A1(_1273_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3026_ (.A1(\beepboop.inst.counter[2] ),
    .A2(_1057_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3027_ (.A1(_0962_),
    .A2(_1058_),
    .A3(_1059_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3028_ (.A1(_1301_),
    .A2(_1057_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3029_ (.A1(_1276_),
    .A2(_1059_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3030_ (.A1(_0962_),
    .A2(_1060_),
    .A3(_1061_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3031_ (.I(_0961_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3032_ (.A1(_1283_),
    .A2(_1059_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3033_ (.A1(_1293_),
    .A2(_1060_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3034_ (.A1(_1062_),
    .A2(_1063_),
    .A3(_1064_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3035_ (.A1(\beepboop.inst.counter[5] ),
    .A2(_1063_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3036_ (.A1(_1291_),
    .A2(_1063_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3037_ (.A1(_1062_),
    .A2(_1065_),
    .A3(_1066_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3038_ (.I(_0961_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3039_ (.A1(_1297_),
    .A2(_1065_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3040_ (.A1(_1067_),
    .A2(_1068_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3041_ (.A1(_1297_),
    .A2(_1065_),
    .B(_1295_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3042_ (.A1(_1284_),
    .A2(\beepboop.inst.counter[6] ),
    .A3(_1065_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3043_ (.A1(_1062_),
    .A2(_1069_),
    .A3(_1070_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3044_ (.A1(_1304_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3045_ (.A1(_1067_),
    .A2(_1071_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3046_ (.A1(_1304_),
    .A2(_1070_),
    .B(_1306_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3047_ (.A1(\beepboop.inst.counter[9] ),
    .A2(\beepboop.inst.counter[8] ),
    .A3(_1070_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3048_ (.A1(_1062_),
    .A2(_1072_),
    .A3(_1073_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3049_ (.A1(_1303_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3050_ (.A1(_1067_),
    .A2(_1074_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3051_ (.A1(_1303_),
    .A2(_1073_),
    .B(\beepboop.inst.counter[11] ),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3052_ (.A1(_1067_),
    .A2(_1075_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3053_ (.D(_0033_),
    .CLK(net90),
    .Q(\ttA_0.data[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3054_ (.D(_0034_),
    .CLK(net108),
    .Q(\ttA_0.data[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3055_ (.D(_0035_),
    .CLK(net103),
    .Q(\ttA_0.data[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3056_ (.D(_0036_),
    .CLK(net108),
    .Q(\ttA_0.data[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3057_ (.D(_0037_),
    .CLK(net103),
    .Q(\ttA_0.data[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3058_ (.D(_0038_),
    .CLK(net108),
    .Q(\ttA_0.data[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3059_ (.D(_0039_),
    .CLK(net103),
    .Q(\ttA_0.data[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3060_ (.D(_0040_),
    .CLK(net108),
    .Q(\ttA_0.data[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3061_ (.D(_0041_),
    .CLK(net68),
    .Q(\ttA_1.top.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3062_ (.D(_0042_),
    .CLK(net68),
    .Q(\ttA_1.top.data[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3063_ (.D(_0043_),
    .CLK(net73),
    .Q(\ttA_1.top.data[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3064_ (.D(_0044_),
    .CLK(net74),
    .Q(\ttA_1.top.data[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3065_ (.D(_0045_),
    .CLK(net73),
    .Q(\ttA_1.top.data[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3066_ (.D(_0046_),
    .CLK(net74),
    .Q(\ttA_1.top.data[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3067_ (.D(_0047_),
    .CLK(net73),
    .Q(\ttA_1.top.data[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3068_ (.D(_0048_),
    .CLK(net69),
    .Q(\ttA_1.top.data[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3069_ (.D(_0049_),
    .CLK(net69),
    .Q(\ttA_1.top.data[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3070_ (.D(_0050_),
    .CLK(net42),
    .Q(\ttA_1.top.data[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3071_ (.D(_0051_),
    .CLK(net42),
    .Q(\ttA_1.top.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3072_ (.D(_0052_),
    .CLK(net43),
    .Q(\ttA_1.top.data[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3073_ (.D(_0053_),
    .CLK(net45),
    .Q(\ttA_1.top.data[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3074_ (.D(_0054_),
    .CLK(net66),
    .Q(\ttA_1.top.data[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3075_ (.D(_0055_),
    .CLK(net45),
    .Q(\ttA_1.top.data[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3076_ (.D(_0056_),
    .CLK(net66),
    .Q(\ttA_1.top.data[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3077_ (.D(_0057_),
    .CLK(net67),
    .Q(\ttA_1.top.data[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3078_ (.D(_0058_),
    .CLK(net66),
    .Q(\ttA_1.top.data[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3079_ (.D(_0059_),
    .CLK(net46),
    .Q(\ttA_1.top.data[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3080_ (.D(_0060_),
    .CLK(net67),
    .Q(\ttA_1.top.data[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3081_ (.D(_0061_),
    .CLK(net46),
    .Q(\ttA_1.top.data[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3082_ (.D(_0062_),
    .CLK(net106),
    .Q(\ttA_0.data[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3083_ (.D(_0063_),
    .CLK(net106),
    .Q(\ttA_0.data[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3084_ (.D(_0064_),
    .CLK(net111),
    .Q(\ttA_0.data[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3085_ (.D(_0065_),
    .CLK(net107),
    .Q(\ttA_0.data[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3086_ (.D(_0066_),
    .CLK(net112),
    .Q(\ttA_0.data[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3087_ (.D(_0067_),
    .CLK(net109),
    .Q(\ttA_0.data[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3088_ (.D(_0068_),
    .CLK(net112),
    .Q(\ttA_0.data[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3089_ (.D(_0069_),
    .CLK(net109),
    .Q(\ttA_0.data[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3090_ (.D(_0070_),
    .CLK(net111),
    .Q(\ttA_0.data[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3091_ (.D(_0071_),
    .CLK(net111),
    .Q(\ttA_0.data[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3092_ (.D(_0072_),
    .CLK(net111),
    .Q(\ttA_0.data[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3093_ (.D(_0073_),
    .CLK(net116),
    .Q(\ttA_0.data[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3094_ (.D(_0074_),
    .CLK(net113),
    .Q(\ttA_0.data[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3095_ (.D(_0075_),
    .CLK(net113),
    .Q(\ttA_0.data[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3096_ (.D(_0076_),
    .CLK(net113),
    .Q(\ttA_0.data[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3097_ (.D(_0077_),
    .CLK(net113),
    .Q(\ttA_0.data[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3098_ (.D(_0078_),
    .CLK(net114),
    .Q(\ttA_0.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3099_ (.D(_0079_),
    .CLK(net114),
    .Q(\ttA_0.data[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3100_ (.D(_0080_),
    .CLK(net114),
    .Q(\ttA_0.data[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3101_ (.D(_0081_),
    .CLK(net115),
    .Q(\ttA_0.data[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3102_ (.D(_0082_),
    .CLK(net112),
    .Q(\ttA_0.data[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3103_ (.D(_0083_),
    .CLK(net112),
    .Q(\ttA_0.data[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3104_ (.D(_0084_),
    .CLK(net115),
    .Q(\ttA_0.data[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3105_ (.D(_0085_),
    .CLK(net110),
    .Q(\ttA_0.data[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3106_ (.D(_0086_),
    .CLK(net83),
    .Q(\ttA_0.prog[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3107_ (.D(_0087_),
    .CLK(net59),
    .Q(\ttA_0.prog[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3108_ (.D(_0088_),
    .CLK(net61),
    .Q(\ttA_0.prog[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3109_ (.D(_0089_),
    .CLK(net84),
    .Q(\ttA_0.prog[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3110_ (.D(_0090_),
    .CLK(net92),
    .Q(\ttA_0.prog[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3111_ (.D(_0091_),
    .CLK(net72),
    .Q(\ttA_0.prog[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3112_ (.D(_0092_),
    .CLK(net71),
    .Q(\ttA_0.prog[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3113_ (.D(_0093_),
    .CLK(net92),
    .Q(\ttA_0.prog[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3114_ (.D(_0094_),
    .CLK(net92),
    .Q(\ttA_0.prog[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3115_ (.D(_0095_),
    .CLK(net72),
    .Q(\ttA_0.prog[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3116_ (.D(_0096_),
    .CLK(net71),
    .Q(\ttA_0.prog[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3117_ (.D(_0097_),
    .CLK(net92),
    .Q(\ttA_0.prog[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3118_ (.D(_0098_),
    .CLK(net71),
    .Q(\ttA_0.prog[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3119_ (.D(_0099_),
    .CLK(net65),
    .Q(\ttA_0.prog[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3120_ (.D(_0100_),
    .CLK(net65),
    .Q(\ttA_0.prog[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3121_ (.D(_0101_),
    .CLK(net71),
    .Q(\ttA_0.prog[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3122_ (.D(_0102_),
    .CLK(net41),
    .Q(\ttA_0.prog[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3123_ (.D(_0103_),
    .CLK(net42),
    .Q(\ttA_0.prog[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3124_ (.D(_0104_),
    .CLK(net41),
    .Q(\ttA_0.prog[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3125_ (.D(_0105_),
    .CLK(net42),
    .Q(\ttA_0.prog[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3126_ (.D(_0106_),
    .CLK(net33),
    .Q(\ttA_0.prog[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3127_ (.D(_0107_),
    .CLK(net64),
    .Q(\ttA_0.prog[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3128_ (.D(_0108_),
    .CLK(net33),
    .Q(\ttA_0.prog[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3129_ (.D(_0109_),
    .CLK(net33),
    .Q(\ttA_0.prog[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3130_ (.D(_0110_),
    .CLK(net41),
    .Q(\ttA_0.prog[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3131_ (.D(_0111_),
    .CLK(net64),
    .Q(\ttA_0.prog[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3132_ (.D(_0112_),
    .CLK(net33),
    .Q(\ttA_0.prog[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3133_ (.D(_0113_),
    .CLK(net36),
    .Q(\ttA_0.prog[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3134_ (.D(_0114_),
    .CLK(net34),
    .Q(\ttA_0.prog[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3135_ (.D(_0115_),
    .CLK(net54),
    .Q(\ttA_0.prog[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3136_ (.D(_0116_),
    .CLK(net35),
    .Q(\ttA_0.prog[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3137_ (.D(_0117_),
    .CLK(net35),
    .Q(\ttA_0.prog[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3138_ (.D(_0118_),
    .CLK(net35),
    .Q(\ttA_0.prog[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3139_ (.D(_0119_),
    .CLK(net54),
    .Q(\ttA_0.prog[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3140_ (.D(_0120_),
    .CLK(net54),
    .Q(\ttA_0.prog[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3141_ (.D(_0121_),
    .CLK(net35),
    .Q(\ttA_0.prog[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3142_ (.D(_0122_),
    .CLK(net60),
    .Q(\ttA_0.prog[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3143_ (.D(_0123_),
    .CLK(net54),
    .Q(\ttA_0.prog[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3144_ (.D(_0124_),
    .CLK(net55),
    .Q(\ttA_0.prog[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3145_ (.D(_0125_),
    .CLK(net60),
    .Q(\ttA_0.prog[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3146_ (.D(_0126_),
    .CLK(net60),
    .Q(\ttA_0.prog[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3147_ (.D(_0127_),
    .CLK(net55),
    .Q(\ttA_0.prog[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3148_ (.D(_0128_),
    .CLK(net55),
    .Q(\ttA_0.prog[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3149_ (.D(_0129_),
    .CLK(net60),
    .Q(\ttA_0.prog[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3150_ (.D(_0130_),
    .CLK(net59),
    .Q(\ttA_0.prog[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3151_ (.D(_0131_),
    .CLK(net59),
    .Q(\ttA_0.prog[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3152_ (.D(_0132_),
    .CLK(net59),
    .Q(\ttA_0.prog[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3153_ (.D(_0133_),
    .CLK(net83),
    .Q(\ttA_0.prog[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3154_ (.D(_0134_),
    .CLK(net95),
    .Q(\ttA_1.top.data[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3155_ (.D(_0135_),
    .CLK(net75),
    .Q(\ttA_1.top.data[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3156_ (.D(_0136_),
    .CLK(net75),
    .Q(\ttA_1.top.data[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3157_ (.D(_0137_),
    .CLK(net109),
    .Q(\ttA_0.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3158_ (.D(_0138_),
    .CLK(net118),
    .Q(\ttA_0.io_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3159_ (.D(_0139_),
    .CLK(net123),
    .Q(\ttA_0.io_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3160_ (.D(_0140_),
    .CLK(net118),
    .Q(\ttA_0.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3161_ (.D(_0141_),
    .CLK(net88),
    .Q(\ttA_0.data[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3162_ (.D(_0142_),
    .CLK(net104),
    .Q(\ttA_0.data[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3163_ (.D(_0143_),
    .CLK(net104),
    .Q(\ttA_0.data[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3164_ (.D(_0144_),
    .CLK(net88),
    .Q(\ttA_0.data[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3165_ (.D(_0145_),
    .RN(_0000_),
    .CLK(net94),
    .Q(\ttA_2.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3166_ (.D(_0146_),
    .RN(_0001_),
    .CLK(net74),
    .Q(\ttA_2.io_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3167_ (.D(_0147_),
    .RN(_0002_),
    .CLK(net73),
    .Q(\ttA_2.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3168_ (.D(_0148_),
    .CLK(net88),
    .Q(\ttA_0.data[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3169_ (.D(_0149_),
    .CLK(net89),
    .Q(\ttA_0.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3170_ (.D(_0150_),
    .CLK(net103),
    .Q(\ttA_0.data[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3171_ (.D(_0151_),
    .CLK(net105),
    .Q(\ttA_0.data[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3172_ (.D(_0152_),
    .CLK(net106),
    .Q(\ttA_0.data[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3173_ (.D(_0153_),
    .CLK(net106),
    .Q(\ttA_0.data[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3174_ (.D(_0154_),
    .CLK(net104),
    .Q(\ttA_0.data[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3175_ (.D(_0155_),
    .CLK(net104),
    .Q(\ttA_0.data[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3176_ (.D(_0156_),
    .CLK(net88),
    .Q(\ttA_0.data[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3177_ (.D(_0157_),
    .CLK(net86),
    .Q(\ttA_0.data[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3178_ (.D(_0158_),
    .CLK(net86),
    .Q(\ttA_0.data[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3179_ (.D(_0159_),
    .CLK(net86),
    .Q(\ttA_0.data[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3180_ (.D(_0160_),
    .CLK(net80),
    .Q(\ttA_0.data[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3181_ (.D(_0161_),
    .CLK(net80),
    .Q(\ttA_0.data[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3182_ (.D(_0162_),
    .CLK(net80),
    .Q(\ttA_0.data[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3183_ (.D(_0163_),
    .CLK(net80),
    .Q(\ttA_0.data[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3184_ (.D(_0164_),
    .CLK(net53),
    .Q(\ttA_0.prog[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3185_ (.D(_0165_),
    .CLK(net53),
    .Q(\ttA_0.prog[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3186_ (.D(_0166_),
    .CLK(net53),
    .Q(\ttA_0.prog[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3187_ (.D(_0167_),
    .CLK(net37),
    .Q(\ttA_0.prog[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3188_ (.D(\ttA_1.top.frontend.rptr_gray1[0] ),
    .RN(_0003_),
    .CLK(net45),
    .Q(\ttA_1.top.frontend.rptr_gray2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3189_ (.D(\ttA_1.top.frontend.rptr_gray1[1] ),
    .RN(_0004_),
    .CLK(net38),
    .Q(\ttA_1.top.frontend.rptr_gray2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3190_ (.D(\ttA_1.top.frontend.rptr_gray1[2] ),
    .RN(_0005_),
    .CLK(net38),
    .Q(\ttA_1.top.frontend.rptr_gray2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3191_ (.D(\ttA_1.top.frontend.rptr_gray1[3] ),
    .RN(_0006_),
    .CLK(net38),
    .Q(\ttA_1.top.frontend.rptr_gray2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3192_ (.D(\ttA_1.top.backend.rptr_b2g.gray[0] ),
    .RN(_0007_),
    .CLK(net47),
    .Q(\ttA_1.top.frontend.rptr_gray1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3193_ (.D(\ttA_1.top.backend.rptr_b2g.gray[1] ),
    .RN(_0008_),
    .CLK(net39),
    .Q(\ttA_1.top.frontend.rptr_gray1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3194_ (.D(\ttA_1.top.backend.rptr_b2g.gray[2] ),
    .RN(_0009_),
    .CLK(net39),
    .Q(\ttA_1.top.frontend.rptr_gray1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3195_ (.D(\ttA_1.top.backend.rptr[3] ),
    .RN(_0010_),
    .CLK(net38),
    .Q(\ttA_1.top.frontend.rptr_gray1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3196_ (.D(_0168_),
    .RN(_0011_),
    .CLK(net30),
    .Q(\ttA_1.top.backend.rptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3197_ (.D(_0169_),
    .RN(_0012_),
    .CLK(net31),
    .Q(\ttA_1.top.backend.rptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3198_ (.D(_0170_),
    .RN(_0013_),
    .CLK(net30),
    .Q(\ttA_1.top.backend.rptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3199_ (.D(_0171_),
    .RN(_0014_),
    .CLK(net31),
    .Q(\ttA_1.top.backend.rptr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3200_ (.D(_0172_),
    .CLK(net81),
    .Q(\ttA_0.data[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3201_ (.D(_0173_),
    .CLK(net83),
    .Q(\ttA_0.data[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3202_ (.D(_0174_),
    .CLK(net82),
    .Q(\ttA_0.data[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3203_ (.D(_0175_),
    .CLK(net84),
    .Q(\ttA_0.data[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3204_ (.D(\ttA_1.top.backend.wptr_gray1[0] ),
    .RN(_0015_),
    .CLK(net31),
    .Q(\ttA_1.top.backend.wptr_gray2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3205_ (.D(\ttA_1.top.backend.wptr_gray1[1] ),
    .RN(_0016_),
    .CLK(net28),
    .Q(\ttA_1.top.backend.wptr_gray2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3206_ (.D(\ttA_1.top.backend.wptr_gray1[2] ),
    .RN(_0017_),
    .CLK(net29),
    .Q(\ttA_1.top.backend.wptr_gray2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3207_ (.D(\ttA_1.top.backend.wptr_gray1[3] ),
    .RN(_0018_),
    .CLK(net29),
    .Q(\ttA_1.top.backend.wptr_gray2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3208_ (.D(\ttA_1.top.backend.wptr_gray[0] ),
    .RN(_0019_),
    .CLK(net29),
    .Q(\ttA_1.top.backend.wptr_gray1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3209_ (.D(\ttA_1.top.backend.wptr_gray[1] ),
    .RN(_0020_),
    .CLK(net28),
    .Q(\ttA_1.top.backend.wptr_gray1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3210_ (.D(\ttA_1.top.backend.wptr_gray[2] ),
    .RN(_0021_),
    .CLK(net28),
    .Q(\ttA_1.top.backend.wptr_gray1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3211_ (.D(\ttA_1.top.backend.wptr_gray[3] ),
    .RN(_0022_),
    .CLK(net28),
    .Q(\ttA_1.top.backend.wptr_gray1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3212_ (.D(_0176_),
    .CLK(net93),
    .Q(\ttA_0.lastdata3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3213_ (.D(net3),
    .RN(_0023_),
    .CLK(net74),
    .Q(\ttA_2.state ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3214_ (.D(_0177_),
    .CLK(net97),
    .Q(\ttA_4.pwm_signal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3215_ (.D(_0178_),
    .CLK(net51),
    .Q(\ttA_0.prog[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3216_ (.D(_0179_),
    .CLK(net51),
    .Q(\ttA_0.prog[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3217_ (.D(_0180_),
    .CLK(net51),
    .Q(\ttA_0.prog[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3218_ (.D(_0181_),
    .CLK(net51),
    .Q(\ttA_0.prog[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3219_ (.D(_0182_),
    .RN(_0024_),
    .CLK(net41),
    .Q(\ttA_1.top.frontend.wptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3220_ (.D(_0183_),
    .RN(_0025_),
    .CLK(net47),
    .Q(\ttA_1.top.frontend.wptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3221_ (.D(_0184_),
    .RN(_0026_),
    .CLK(net45),
    .Q(\ttA_1.top.frontend.wptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3222_ (.D(_0185_),
    .RN(_0027_),
    .CLK(net44),
    .Q(\ttA_1.top.backend.wptr_gray[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3223_ (.D(_0186_),
    .CLK(net97),
    .Q(\ttA_6.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3224_ (.D(_0187_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3225_ (.D(_0188_),
    .CLK(net57),
    .Q(\ttA_0.prog[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3226_ (.D(_0189_),
    .CLK(net57),
    .Q(\ttA_0.prog[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3227_ (.D(_0190_),
    .CLK(net52),
    .Q(\ttA_0.prog[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3228_ (.D(_0191_),
    .CLK(net57),
    .Q(\ttA_0.prog[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3229_ (.D(_0192_),
    .CLK(net58),
    .Q(\ttA_0.prog[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3230_ (.D(_0193_),
    .CLK(net58),
    .Q(\ttA_0.prog[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3231_ (.D(_0194_),
    .CLK(net57),
    .Q(\ttA_0.prog[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3232_ (.D(_0195_),
    .CLK(net58),
    .Q(\ttA_0.prog[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3233_ (.D(_0196_),
    .CLK(net118),
    .Q(\ttA_4.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3234_ (.D(_0197_),
    .CLK(net118),
    .Q(\ttA_4.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3235_ (.D(_0198_),
    .CLK(net122),
    .Q(\ttA_4.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3236_ (.D(_0199_),
    .CLK(net121),
    .Q(\ttA_4.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3237_ (.D(_0200_),
    .CLK(net119),
    .Q(\ttA_4.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3238_ (.D(_0201_),
    .CLK(net119),
    .Q(\ttA_4.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3239_ (.D(_0202_),
    .CLK(net82),
    .Q(\ttA_0.data[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3240_ (.D(_0203_),
    .CLK(net81),
    .Q(\ttA_0.data[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3241_ (.D(_0204_),
    .CLK(net82),
    .Q(\ttA_0.data[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3242_ (.D(_0205_),
    .CLK(net85),
    .Q(\ttA_0.data[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3243_ (.D(_0206_),
    .CLK(net97),
    .Q(\ttA_4.active_duty[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3244_ (.D(_0207_),
    .CLK(net94),
    .Q(\ttA_4.active_duty[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3245_ (.D(_0208_),
    .CLK(net100),
    .Q(\ttA_4.active_duty[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3246_ (.D(_0209_),
    .CLK(net99),
    .Q(\ttA_4.active_duty[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3247_ (.D(_0210_),
    .CLK(net100),
    .Q(\ttA_4.active_duty[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3248_ (.D(_0211_),
    .CLK(net97),
    .Q(\ttA_4.active_duty[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3249_ (.D(_0212_),
    .CLK(net83),
    .Q(\ttA_0.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3250_ (.D(_0213_),
    .CLK(net93),
    .Q(\ttA_0.io_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3251_ (.D(_0214_),
    .CLK(net93),
    .Q(\ttA_0.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3252_ (.D(_0215_),
    .CLK(net93),
    .Q(\ttA_0.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3253_ (.D(_0216_),
    .CLK(net86),
    .Q(\ttA_0.data[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3254_ (.D(_0217_),
    .CLK(net87),
    .Q(\ttA_0.data[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3255_ (.D(_0218_),
    .CLK(net87),
    .Q(\ttA_0.data[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3256_ (.D(_0219_),
    .CLK(net90),
    .Q(\ttA_0.data[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3257_ (.D(_0220_),
    .CLK(net99),
    .Q(\ttA_6.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3258_ (.D(_0221_),
    .CLK(net121),
    .Q(\ttA_6.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3259_ (.D(_0222_),
    .CLK(net119),
    .Q(\ttA_6.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3260_ (.D(_0223_),
    .CLK(net119),
    .Q(\ttA_6.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3261_ (.D(_0224_),
    .CLK(net120),
    .Q(\ttA_6.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3262_ (.D(_0225_),
    .CLK(net120),
    .Q(\ttA_6.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3263_ (.D(_0226_),
    .CLK(net121),
    .Q(\ttA_6.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3264_ (.D(_0227_),
    .CLK(net100),
    .Q(\ttA_6.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3265_ (.D(_0228_),
    .CLK(net98),
    .Q(\ttA_6.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3266_ (.D(_0229_),
    .CLK(net98),
    .Q(\ttA_6.counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3267_ (.D(_0230_),
    .CLK(net96),
    .Q(\ttA_6.counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3268_ (.D(net294),
    .CLK(net123),
    .Q(\ttA_6.counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3269_ (.D(net293),
    .CLK(net123),
    .Q(\ttA_6.counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3270_ (.D(net292),
    .CLK(net123),
    .Q(\ttA_6.counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3271_ (.D(net291),
    .CLK(net124),
    .Q(\ttA_6.counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3272_ (.D(_0235_),
    .RN(_0028_),
    .CLK(net66),
    .Q(\ttA_2.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3273_ (.D(_0236_),
    .RN(_0029_),
    .CLK(net64),
    .Q(\ttA_2.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3274_ (.D(_0237_),
    .RN(_0030_),
    .CLK(net43),
    .Q(\ttA_2.io_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3275_ (.D(_0238_),
    .RN(_0031_),
    .CLK(net64),
    .Q(\ttA_2.io_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _3276_ (.D(_0239_),
    .RN(_0032_),
    .CLK(net65),
    .Q(\ttA_2.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3277_ (.D(_0240_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3278_ (.D(_0241_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3279_ (.D(_0242_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3280_ (.D(_0243_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3281_ (.D(_0244_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3282_ (.D(_0245_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3283_ (.D(_0246_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3284_ (.D(_0247_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3285_ (.D(_0248_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3286_ (.D(_0249_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3287_ (.D(_0250_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3288_ (.D(net290),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3289_ (.D(net289),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3290_ (.D(net288),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3291_ (.D(net287),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\beepboop.inst.counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_296 (.Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_297 (.Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_236 (.ZN(net236));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_237 (.ZN(net237));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_238 (.ZN(net238));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_239 (.ZN(net239));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_240 (.ZN(net240));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_241 (.ZN(net241));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_242 (.ZN(net242));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_243 (.ZN(net243));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_244 (.ZN(net244));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_245 (.ZN(net245));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_246 (.ZN(net246));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_247 (.ZN(net247));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_248 (.ZN(net248));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_249 (.ZN(net249));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_250 (.ZN(net250));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_251 (.ZN(net251));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_252 (.ZN(net252));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_253 (.ZN(net253));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_254 (.ZN(net254));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_255 (.ZN(net255));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_256 (.ZN(net256));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_257 (.ZN(net257));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_258 (.ZN(net258));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_259 (.ZN(net259));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_260 (.ZN(net260));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_261 (.ZN(net261));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_262 (.ZN(net262));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_263 (.ZN(net263));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_264 (.ZN(net264));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_265 (.ZN(net265));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_266 (.ZN(net266));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_267 (.ZN(net267));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_268 (.ZN(net268));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_269 (.ZN(net269));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_270 (.ZN(net270));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_271 (.ZN(net271));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_272 (.ZN(net272));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_273 (.ZN(net273));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_274 (.ZN(net274));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_275 (.ZN(net275));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_276 (.ZN(net276));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_277 (.ZN(net277));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_278 (.ZN(net278));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_279 (.ZN(net279));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_280 (.ZN(net280));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_281 (.ZN(net281));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_282 (.ZN(net282));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_283 (.ZN(net283));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_284 (.ZN(net284));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_285 (.ZN(net285));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_286 (.ZN(net286));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3291__287 (.ZN(net287));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3290__288 (.ZN(net288));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3289__289 (.ZN(net289));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3288__290 (.ZN(net290));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3271__291 (.ZN(net291));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3270__292 (.ZN(net292));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3269__293 (.ZN(net293));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3268__294 (.ZN(net294));
 gf180mcu_fd_sc_mcu7t5v0__tieh user_proj_295 (.Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3462_ (.I(net27),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input5 (.I(io_in[14]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[15]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input8 (.I(io_in[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_in[20]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_in[30]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(io_in[31]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout28 (.I(net30),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout29 (.I(net30),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout32 (.I(net2),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(net36),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout36 (.I(net37),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout37 (.I(net50),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net40),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout40 (.I(net49),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net44),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout42 (.I(net44),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(net44),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(net48),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net47),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout46 (.I(net47),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net79),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net56),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout54 (.I(net56),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net63),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net62),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net62),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net62),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net63),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout63 (.I(net78),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout64 (.I(net70),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net70),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout66 (.I(net68),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net70),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net77),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout71 (.I(net76),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net76),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout73 (.I(net75),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net76),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net79),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout79 (.I(net127),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net81),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout82 (.I(net85),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout85 (.I(net91),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout86 (.I(net89),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net89),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout90 (.I(net91),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout91 (.I(net102),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout92 (.I(net94),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net96),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net96),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net101),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net99),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net101),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout101 (.I(net102),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net126),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net105),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net107),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout105 (.I(net107),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net110),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout109 (.I(net110),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout110 (.I(net117),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout111 (.I(net116),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net115),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout113 (.I(net114),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net116),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net125),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net122),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout119 (.I(net122),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout120 (.I(net121),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout121 (.I(net122),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout122 (.I(net124),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net125),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout125 (.I(net126),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net127),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net1),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel user_proj_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__RN (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A2 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A2 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__B (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__RN (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A1 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__D (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__D (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__D (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__D (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__I (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__C (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A1 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A1 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__S0 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__I (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__S0 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__S0 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__S0 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A2 (.I(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__S0 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__S0 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__S0 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__S0 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2081__I (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__I (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2041__I (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__I (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__S0 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__S1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__S1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__S1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__I (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__S0 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__I (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__S1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__S1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2023__A2 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A2 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2027__A2 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A3 (.I(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2033__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2065__I (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__B (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__B (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2037__B (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__S1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__S1 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__S0 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__S0 (.I(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__S1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__S1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__S1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__S1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__S0 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__S0 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__S0 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__S0 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__S1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__S1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__S1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__S1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__B (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A2 (.I(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__S0 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__S0 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__S0 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__S0 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__S0 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__S1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__S0 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__S1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__S1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__S1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__S0 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__S0 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__S1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__S1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__S1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__S1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__B (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__I (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__I (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__I (.I(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__B (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__C (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__I (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__I (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__C (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__C (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__C (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A3 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__I (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__I (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__I (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2158__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__I (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__C (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__I (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__B2 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__A1 (.I(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__I (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__A1 (.I(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__I (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__A3 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A3 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__C (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__C (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__C (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__C (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__I (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__C (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__C (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__C (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__C (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__I (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A2 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__C (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__C (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__C (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__B2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__I (.I(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__I (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__B (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__B (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__I (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2866__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__B (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__B (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2887__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2860__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__B (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A3 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A3 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__B1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__C (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__C (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__B (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A4 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A3 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__C (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__B1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A2 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A3 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__I (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__B (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__B (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__B (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A3 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A3 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__B (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__B (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A3 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__C (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__B (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__B1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__B2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__B (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__B1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__C (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__C (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A2 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__C (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A3 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__B (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__C (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A3 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3017__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__C (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__C (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__C (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__C (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2979__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2983__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__I (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2807__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__I (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2810__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2808__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__I (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__I (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__I (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__B (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2834__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__B1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__A3 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__B2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A2 (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__I (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__B (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A2 (.I(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__B (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__B (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__B (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__B (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__A4 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__I (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__I (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2947__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__B (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__A3 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2987__I (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__A3 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A3 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3048__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3043__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3052__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3050__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__B (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__B2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A3 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A2 (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__I (.I(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__I (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__B1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__B2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__B (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__C (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__B2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A3 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__B2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__I1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__B2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1629__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A2 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__B (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__C (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A3 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__I (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__I (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__B (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__B (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A3 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__B (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A3 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__B1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__I (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__I (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__B (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__C (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__I (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A3 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__C (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__C (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__I0 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A4 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A3 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__B (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__B (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A3 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A4 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1798__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__S0 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__S0 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__I (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__I (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__S0 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__S0 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__S0 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__I (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__S1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__S1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__S0 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__I (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__C2 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__I (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__C (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__I (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__I (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__I (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__I (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__B2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2993__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A1 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__C (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A2 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A3 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A3 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__S1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__S1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__S1 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__I (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__S1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__S1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__S1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__I (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__S0 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__S0 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__S1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__I (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__B (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__A2 (.I(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__I (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1884__B1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2093__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__B2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__B2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__B (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__C (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__I (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2067__B (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__B2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__B (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__C (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A3 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A4 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__B2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__B2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__S0 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A1 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__S0 (.I(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__S1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__S1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__C (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__S1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__S0 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__S (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__B (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__B (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__I (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2152__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__B (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(\ttA_0.data[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__I0 (.I(\ttA_0.data[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__A1 (.I(\ttA_0.data[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I0 (.I(\ttA_0.data[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(\ttA_0.data[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__I0 (.I(\ttA_0.data[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A1 (.I(\ttA_0.data[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__I2 (.I(\ttA_0.data[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(\ttA_0.data[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I2 (.I(\ttA_0.data[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(\ttA_0.data[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I2 (.I(\ttA_0.data[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__A1 (.I(\ttA_0.data[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I2 (.I(\ttA_0.data[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(\ttA_0.data[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__I0 (.I(\ttA_0.data[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__A1 (.I(\ttA_0.data[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__I0 (.I(\ttA_0.data[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(\ttA_0.data[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I0 (.I(\ttA_0.data[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(\ttA_0.data[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__I0 (.I(\ttA_0.data[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__A1 (.I(\ttA_0.data[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__I2 (.I(\ttA_0.data[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__A1 (.I(\ttA_0.data[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__I2 (.I(\ttA_0.data[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A1 (.I(\ttA_0.data[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__I1 (.I(\ttA_0.data[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(\ttA_0.data[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__I1 (.I(\ttA_0.data[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(\ttA_0.data[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__I1 (.I(\ttA_0.data[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A1 (.I(\ttA_0.data[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I1 (.I(\ttA_0.data[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2814__A1 (.I(\ttA_0.data[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__I2 (.I(\ttA_0.data[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(\ttA_0.data[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I2 (.I(\ttA_0.data[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2818__A1 (.I(\ttA_0.data[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__I2 (.I(\ttA_0.data[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A1 (.I(\ttA_0.data[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I2 (.I(\ttA_0.data[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A1 (.I(\ttA_0.data[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__I3 (.I(\ttA_0.data[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(\ttA_0.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__I3 (.I(\ttA_0.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(\ttA_0.data[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I3 (.I(\ttA_0.data[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A1 (.I(\ttA_0.data[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__I2 (.I(\ttA_0.data[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(\ttA_0.data[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__I2 (.I(\ttA_0.data[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(\ttA_0.data[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__I2 (.I(\ttA_0.data[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__A1 (.I(\ttA_0.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__I1 (.I(\ttA_0.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(\ttA_0.data[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__I1 (.I(\ttA_0.data[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(\ttA_0.data[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__I1 (.I(\ttA_0.data[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(\ttA_0.data[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__I1 (.I(\ttA_0.data[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(\ttA_0.data[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__I0 (.I(\ttA_0.data[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A1 (.I(\ttA_0.data[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I0 (.I(\ttA_0.data[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(\ttA_0.data[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I0 (.I(\ttA_0.data[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__A1 (.I(\ttA_0.data[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I0 (.I(\ttA_0.data[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__A1 (.I(\ttA_0.data[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__I1 (.I(\ttA_0.data[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(\ttA_0.data[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2112__I1 (.I(\ttA_0.data[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(\ttA_0.data[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I1 (.I(\ttA_0.data[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(\ttA_0.data[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__I1 (.I(\ttA_0.data[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__I (.I(\ttA_0.io_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__I (.I(\ttA_0.io_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__I (.I(\ttA_0.io_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__I (.I(\ttA_0.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(\ttA_0.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__I (.I(\ttA_0.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__I (.I(\ttA_0.io_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__I (.I(\ttA_0.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__I (.I(\ttA_0.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__I (.I(\ttA_0.prog[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__I2 (.I(\ttA_0.prog[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__I (.I(\ttA_0.prog[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__I3 (.I(\ttA_0.prog[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__I (.I(\ttA_0.prog[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__I3 (.I(\ttA_0.prog[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(\ttA_0.prog[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__I0 (.I(\ttA_0.prog[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(\ttA_0.prog[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__I0 (.I(\ttA_0.prog[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A1 (.I(\ttA_0.prog[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__I0 (.I(\ttA_0.prog[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(\ttA_0.prog[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__I0 (.I(\ttA_0.prog[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A1 (.I(\ttA_0.prog[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__I1 (.I(\ttA_0.prog[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(\ttA_0.prog[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__I2 (.I(\ttA_0.prog[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__I (.I(\ttA_0.prog[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__I2 (.I(\ttA_0.prog[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__I (.I(\ttA_0.prog[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__I2 (.I(\ttA_0.prog[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__I (.I(\ttA_0.prog[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__I2 (.I(\ttA_0.prog[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__I (.I(\ttA_0.prog[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__I3 (.I(\ttA_0.prog[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__I (.I(\ttA_0.prog[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__I3 (.I(\ttA_0.prog[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__I (.I(\ttA_0.prog[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__I3 (.I(\ttA_0.prog[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__I (.I(\ttA_0.prog[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__I3 (.I(\ttA_0.prog[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(\ttA_0.prog[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__I0 (.I(\ttA_0.prog[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A1 (.I(\ttA_0.prog[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__I0 (.I(\ttA_0.prog[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__I (.I(\ttA_0.prog[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__I3 (.I(\ttA_0.prog[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__I (.I(\ttA_0.prog[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__I3 (.I(\ttA_0.prog[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__C (.I(\ttA_1.top.backend.rptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A1 (.I(\ttA_1.top.backend.rptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1693__A1 (.I(\ttA_1.top.backend.rptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__I (.I(\ttA_1.top.backend.rptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__D (.I(\ttA_1.top.backend.rptr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(\ttA_1.top.backend.rptr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(\ttA_1.top.backend.rptr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__D (.I(\ttA_1.top.backend.rptr_b2g.gray[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(\ttA_1.top.backend.rptr_b2g.gray[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__D (.I(\ttA_1.top.backend.wptr_gray[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(\ttA_1.top.backend.wptr_gray[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(\ttA_1.top.backend.wptr_gray[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__D (.I(\ttA_1.top.backend.wptr_gray[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(\ttA_1.top.backend.wptr_gray[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A1 (.I(\ttA_1.top.backend.wptr_gray[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A1 (.I(\ttA_1.top.backend.wptr_gray[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A1 (.I(\ttA_1.top.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__I1 (.I(\ttA_1.top.data[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(\ttA_1.top.data[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__I0 (.I(\ttA_1.top.data[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__A1 (.I(\ttA_1.top.data[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__I0 (.I(\ttA_1.top.data[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A1 (.I(\ttA_1.top.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__I2 (.I(\ttA_1.top.data[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A1 (.I(\ttA_1.top.data[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__I3 (.I(\ttA_1.top.data[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(\ttA_1.top.frontend.rptr_gray2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A2 (.I(\ttA_1.top.frontend.wptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1686__A1 (.I(\ttA_1.top.frontend.wptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(\ttA_1.top.frontend.wptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A2 (.I(\ttA_1.top.frontend.wptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__I (.I(\ttA_1.top.frontend.wptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(\ttA_1.top.frontend.wptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A2 (.I(\ttA_1.top.frontend.wptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__I (.I(\ttA_1.top.frontend.wptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__I (.I(\ttA_1.top.frontend.wptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(\ttA_1.top.frontend.wptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1660__A2 (.I(\ttA_1.top.frontend.wptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__I (.I(\ttA_1.top.frontend.wptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__B2 (.I(\ttA_2.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I (.I(\ttA_2.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A2 (.I(\ttA_2.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A2 (.I(\ttA_2.io_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A1 (.I(\ttA_2.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(\ttA_2.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A1 (.I(\ttA_2.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__I (.I(\ttA_2.io_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(\ttA_2.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__I (.I(\ttA_2.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A1 (.I(\ttA_2.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A1 (.I(\ttA_2.io_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A1 (.I(\ttA_2.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__A1 (.I(\ttA_2.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__A1 (.I(\ttA_2.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A1 (.I(\ttA_2.io_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2946__A1 (.I(\ttA_4.active_duty[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__B (.I(\ttA_4.active_duty[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__A1 (.I(\ttA_4.active_duty[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__B1 (.I(\ttA_4.active_duty[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(\ttA_4.active_duty[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A1 (.I(\ttA_4.active_duty[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2839__I (.I(\ttA_4.active_duty[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(\ttA_4.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A2 (.I(\ttA_4.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__B2 (.I(\ttA_4.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__I (.I(\ttA_4.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(\ttA_4.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__A1 (.I(\ttA_4.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2854__B2 (.I(\ttA_4.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(\ttA_4.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(\ttA_4.pwm_signal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A1 (.I(\ttA_4.pwm_signal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A1 (.I(\ttA_6.counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(\ttA_6.counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__I (.I(\ttA_6.counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(\ttA_6.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__I (.I(\ttA_6.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(\ttA_6.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__A1 (.I(\ttA_6.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A1 (.I(\ttA_6.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__I (.I(\ttA_6.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__I (.I(\ttA_6.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__D (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__B2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__B (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__B1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__B2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__CLK (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__CLK (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__CLK (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3133__CLK (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3130__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__CLK (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3071__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3070__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__CLK (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__CLK (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__CLK (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3225__CLK (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3107__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__CLK (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__CLK (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__CLK (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__CLK (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3142__CLK (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3076__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__CLK (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3061__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__CLK (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3065__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3063__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__CLK (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3240__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__CLK (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3109__CLK (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__CLK (.I(net86));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3176__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__CLK (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__CLK (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__CLK (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__CLK (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3247__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3059__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3057__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__CLK (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__CLK (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__CLK (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__CLK (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__CLK (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__CLK (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__CLK (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3105__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__CLK (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3235__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[0] = net128;
 assign io_oeb[10] = net295;
 assign io_oeb[11] = net138;
 assign io_oeb[12] = net139;
 assign io_oeb[13] = net140;
 assign io_oeb[14] = net141;
 assign io_oeb[15] = net142;
 assign io_oeb[16] = net143;
 assign io_oeb[17] = net144;
 assign io_oeb[18] = net296;
 assign io_oeb[19] = net145;
 assign io_oeb[1] = net129;
 assign io_oeb[20] = net146;
 assign io_oeb[21] = net147;
 assign io_oeb[22] = net148;
 assign io_oeb[23] = net149;
 assign io_oeb[24] = net150;
 assign io_oeb[25] = net151;
 assign io_oeb[26] = net152;
 assign io_oeb[27] = net153;
 assign io_oeb[28] = net154;
 assign io_oeb[29] = net155;
 assign io_oeb[2] = net130;
 assign io_oeb[30] = net297;
 assign io_oeb[31] = net156;
 assign io_oeb[32] = net157;
 assign io_oeb[33] = net158;
 assign io_oeb[34] = net159;
 assign io_oeb[35] = net160;
 assign io_oeb[36] = net161;
 assign io_oeb[37] = net162;
 assign io_oeb[3] = net131;
 assign io_oeb[4] = net132;
 assign io_oeb[5] = net133;
 assign io_oeb[6] = net134;
 assign io_oeb[7] = net135;
 assign io_oeb[8] = net136;
 assign io_oeb[9] = net137;
 assign io_out[0] = net163;
 assign io_out[10] = net173;
 assign io_out[11] = net174;
 assign io_out[12] = net175;
 assign io_out[13] = net176;
 assign io_out[14] = net177;
 assign io_out[15] = net178;
 assign io_out[16] = net179;
 assign io_out[17] = net180;
 assign io_out[18] = net181;
 assign io_out[19] = net182;
 assign io_out[1] = net164;
 assign io_out[20] = net183;
 assign io_out[29] = net184;
 assign io_out[2] = net165;
 assign io_out[30] = net185;
 assign io_out[31] = net186;
 assign io_out[3] = net166;
 assign io_out[4] = net167;
 assign io_out[5] = net168;
 assign io_out[6] = net169;
 assign io_out[7] = net170;
 assign io_out[8] = net171;
 assign io_out[9] = net172;
 assign irq[0] = net187;
 assign irq[1] = net188;
 assign irq[2] = net189;
 assign la_data_out[0] = net190;
 assign la_data_out[10] = net200;
 assign la_data_out[11] = net201;
 assign la_data_out[12] = net202;
 assign la_data_out[13] = net203;
 assign la_data_out[14] = net204;
 assign la_data_out[15] = net205;
 assign la_data_out[16] = net206;
 assign la_data_out[17] = net207;
 assign la_data_out[18] = net208;
 assign la_data_out[19] = net209;
 assign la_data_out[1] = net191;
 assign la_data_out[20] = net210;
 assign la_data_out[21] = net211;
 assign la_data_out[22] = net212;
 assign la_data_out[23] = net213;
 assign la_data_out[24] = net214;
 assign la_data_out[25] = net215;
 assign la_data_out[26] = net216;
 assign la_data_out[27] = net217;
 assign la_data_out[28] = net218;
 assign la_data_out[29] = net219;
 assign la_data_out[2] = net192;
 assign la_data_out[30] = net220;
 assign la_data_out[31] = net221;
 assign la_data_out[32] = net222;
 assign la_data_out[33] = net223;
 assign la_data_out[34] = net224;
 assign la_data_out[35] = net225;
 assign la_data_out[36] = net226;
 assign la_data_out[37] = net227;
 assign la_data_out[38] = net228;
 assign la_data_out[39] = net229;
 assign la_data_out[3] = net193;
 assign la_data_out[40] = net230;
 assign la_data_out[41] = net231;
 assign la_data_out[42] = net232;
 assign la_data_out[43] = net233;
 assign la_data_out[44] = net234;
 assign la_data_out[45] = net235;
 assign la_data_out[46] = net236;
 assign la_data_out[47] = net237;
 assign la_data_out[48] = net238;
 assign la_data_out[49] = net239;
 assign la_data_out[4] = net194;
 assign la_data_out[50] = net240;
 assign la_data_out[51] = net241;
 assign la_data_out[52] = net242;
 assign la_data_out[53] = net243;
 assign la_data_out[54] = net244;
 assign la_data_out[55] = net245;
 assign la_data_out[56] = net246;
 assign la_data_out[57] = net247;
 assign la_data_out[58] = net248;
 assign la_data_out[59] = net249;
 assign la_data_out[5] = net195;
 assign la_data_out[60] = net250;
 assign la_data_out[61] = net251;
 assign la_data_out[62] = net252;
 assign la_data_out[63] = net253;
 assign la_data_out[6] = net196;
 assign la_data_out[7] = net197;
 assign la_data_out[8] = net198;
 assign la_data_out[9] = net199;
 assign wbs_ack_o = net254;
 assign wbs_dat_o[0] = net255;
 assign wbs_dat_o[10] = net265;
 assign wbs_dat_o[11] = net266;
 assign wbs_dat_o[12] = net267;
 assign wbs_dat_o[13] = net268;
 assign wbs_dat_o[14] = net269;
 assign wbs_dat_o[15] = net270;
 assign wbs_dat_o[16] = net271;
 assign wbs_dat_o[17] = net272;
 assign wbs_dat_o[18] = net273;
 assign wbs_dat_o[19] = net274;
 assign wbs_dat_o[1] = net256;
 assign wbs_dat_o[20] = net275;
 assign wbs_dat_o[21] = net276;
 assign wbs_dat_o[22] = net277;
 assign wbs_dat_o[23] = net278;
 assign wbs_dat_o[24] = net279;
 assign wbs_dat_o[25] = net280;
 assign wbs_dat_o[26] = net281;
 assign wbs_dat_o[27] = net282;
 assign wbs_dat_o[28] = net283;
 assign wbs_dat_o[29] = net284;
 assign wbs_dat_o[2] = net257;
 assign wbs_dat_o[30] = net285;
 assign wbs_dat_o[31] = net286;
 assign wbs_dat_o[3] = net258;
 assign wbs_dat_o[4] = net259;
 assign wbs_dat_o[5] = net260;
 assign wbs_dat_o[6] = net261;
 assign wbs_dat_o[7] = net262;
 assign wbs_dat_o[8] = net263;
 assign wbs_dat_o[9] = net264;
endmodule

